module SYS_TOP
(
 input REF_CLK ,
 input UART_CLK,
 input RST     ,
 input RX_IN   ,

 output TX_OUT
);





///////////////////////////////////////////////////////
///////////////////////////////////////////////////////
//////////////// BLOCKS CONNECTION ////////////////////
///////////////////////////////////////////////////////
///////////////////////////////////////////////////////

endmodule