module SYS_TOP (
	SI, 
	SE, 
	scan_clk, 
	scan_rst, 
	test_mode, 
	SO, 
	REF_CLK, 
	UART_CLK, 
	RST, 
	RX_IN, 
	TX_OUT, 
	test_si2, 
	test_so2, 
	test_si3, 
	test_so3, 
	test_si4, 
	test_so4, 
	test_si5, 
	test_so5);
   input SI;
   input SE;
   input scan_clk;
   input scan_rst;
   input test_mode;
   output SO;
   input REF_CLK;
   input UART_CLK;
   input RST;
   input RX_IN;
   output TX_OUT;
   input test_si2;
   output test_so2;
   input test_si3;
   output test_so3;
   input test_si4;
   output test_so4;
   input test_si5;
   output test_so5;

   // Internal wires
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N1;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N2;
   wire scan_clk__L2_N1;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire REF_CLK_M__L5_N7;
   wire REF_CLK_M__L5_N6;
   wire REF_CLK_M__L5_N5;
   wire REF_CLK_M__L5_N4;
   wire REF_CLK_M__L5_N3;
   wire REF_CLK_M__L5_N2;
   wire REF_CLK_M__L5_N1;
   wire REF_CLK_M__L5_N0;
   wire REF_CLK_M__L4_N0;
   wire REF_CLK_M__L3_N0;
   wire REF_CLK_M__L2_N1;
   wire REF_CLK_M__L2_N0;
   wire REF_CLK_M__L1_N0;
   wire ALU_CLK__L1_N0;
   wire UART_CLK_M__L8_N3;
   wire UART_CLK_M__L8_N2;
   wire UART_CLK_M__L8_N1;
   wire UART_CLK_M__L8_N0;
   wire UART_CLK_M__L7_N0;
   wire UART_CLK_M__L6_N0;
   wire UART_CLK_M__L5_N0;
   wire UART_CLK_M__L4_N0;
   wire UART_CLK_M__L3_N0;
   wire UART_CLK_M__L2_N2;
   wire UART_CLK_M__L2_N1;
   wire UART_CLK_M__L2_N0;
   wire UART_CLK_M__L1_N0;
   wire RX_CLK_M__L1_N0;
   wire TX_CLK_M__L1_N0;
   wire FE_OFN24_SE;
   wire FE_OFN22_SE;
   wire FE_OFN21_SE;
   wire FE_OFN20_SE;
   wire FE_OFN19_SE;
   wire FE_OFN18_SE;
   wire FE_OFN17_SE;
   wire FE_OFN15_RST_D2_M;
   wire FE_OFN14_RST_D2_M;
   wire FE_OFN12_RST_D1_M;
   wire FE_OFN11_RST_D1_M;
   wire FE_OFN10_RST_D1_M;
   wire FE_OFN8_RST_D1_M;
   wire REF_CLK_M;
   wire UART_CLK_M;
   wire RST_M;
   wire RX_CLK;
   wire RX_CLK_M;
   wire TX_CLK;
   wire TX_CLK_M;
   wire RST_D1;
   wire RST_D1_M;
   wire RST_D2;
   wire RST_D2_M;
   wire Gate_En;
   wire ALU_CLK;
   wire in_Data_Sys_en;
   wire enable_pulse;
   wire F_Full;
   wire Rd_Valid;
   wire OUT_VALID;
   wire WR_INC;
   wire Enable;
   wire RdEn;
   wire WrEn;
   wire F_Empty;
   wire busy;
   wire R_INC;
   wire n1;
   wire n2;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n16;
   wire n19;
   wire n20;
   wire n21;
   wire [7:0] REG3;
   wire [7:0] in_Data_Sys;
   wire [7:0] SYNC_bus;
   wire [7:0] RdData;
   wire [15:0] ALU_OUT;
   wire [7:0] WR_DATA;
   wire [3:0] ALU_FUN;
   wire [7:0] Wr_D;
   wire [7:0] Addr;
   wire [7:0] REG0;
   wire [7:0] REG1;
   wire [7:0] REG2;
   wire [7:0] in_DATA_tx;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;
   wire SYNOPSYS_UNCONNECTED__2;
   wire SYNOPSYS_UNCONNECTED__3;

   assign test_so5 = R_INC ;

   CLKINVX40M REF_CLK__L2_I0 (.Y(REF_CLK__L2_N0), 
	.A(REF_CLK__L1_N0));
   CLKINVX40M REF_CLK__L1_I0 (.Y(REF_CLK__L1_N0), 
	.A(REF_CLK));
   CLKINVX40M UART_CLK__L2_I0 (.Y(UART_CLK__L2_N0), 
	.A(UART_CLK__L1_N0));
   CLKINVX40M UART_CLK__L1_I0 (.Y(UART_CLK__L1_N0), 
	.A(UART_CLK));
   INVX2M scan_clk__L5_I0 (.Y(scan_clk__L5_N0), 
	.A(scan_clk__L4_N0));
   CLKINVX1M scan_clk__L4_I0 (.Y(scan_clk__L4_N0), 
	.A(scan_clk__L3_N1));
   CLKINVX1M scan_clk__L3_I1 (.Y(scan_clk__L3_N1), 
	.A(scan_clk__L2_N2));
   INVX2M scan_clk__L3_I0 (.Y(scan_clk__L3_N0), 
	.A(scan_clk__L2_N1));
   CLKBUFX3M scan_clk__L2_I2 (.Y(scan_clk__L2_N2), 
	.A(scan_clk__L1_N0));
   BUFX3M scan_clk__L2_I1 (.Y(scan_clk__L2_N1), 
	.A(scan_clk__L1_N0));
   INVX2M scan_clk__L2_I0 (.Y(scan_clk__L2_N0), 
	.A(scan_clk__L1_N0));
   CLKINVX40M scan_clk__L1_I0 (.Y(scan_clk__L1_N0), 
	.A(scan_clk));
   CLKINVX12M REF_CLK_M__L5_I7 (.Y(REF_CLK_M__L5_N7), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX12M REF_CLK_M__L5_I6 (.Y(REF_CLK_M__L5_N6), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX12M REF_CLK_M__L5_I5 (.Y(REF_CLK_M__L5_N5), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX12M REF_CLK_M__L5_I4 (.Y(REF_CLK_M__L5_N4), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX12M REF_CLK_M__L5_I3 (.Y(REF_CLK_M__L5_N3), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX12M REF_CLK_M__L5_I2 (.Y(REF_CLK_M__L5_N2), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX12M REF_CLK_M__L5_I1 (.Y(REF_CLK_M__L5_N1), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX12M REF_CLK_M__L5_I0 (.Y(REF_CLK_M__L5_N0), 
	.A(REF_CLK_M__L4_N0));
   CLKINVX32M REF_CLK_M__L4_I0 (.Y(REF_CLK_M__L4_N0), 
	.A(REF_CLK_M__L3_N0));
   CLKINVX40M REF_CLK_M__L3_I0 (.Y(REF_CLK_M__L3_N0), 
	.A(REF_CLK_M__L2_N1));
   CLKBUFX40M REF_CLK_M__L2_I1 (.Y(REF_CLK_M__L2_N1), 
	.A(REF_CLK_M__L1_N0));
   CLKINVX12M REF_CLK_M__L2_I0 (.Y(REF_CLK_M__L2_N0), 
	.A(REF_CLK_M__L1_N0));
   CLKINVX3M REF_CLK_M__L1_I0 (.Y(REF_CLK_M__L1_N0), 
	.A(REF_CLK_M));
   CLKBUFX40M ALU_CLK__L1_I0 (.Y(ALU_CLK__L1_N0), 
	.A(ALU_CLK));
   INVX6M UART_CLK_M__L8_I3 (.Y(UART_CLK_M__L8_N3), 
	.A(UART_CLK_M__L7_N0));
   INVX6M UART_CLK_M__L8_I2 (.Y(UART_CLK_M__L8_N2), 
	.A(UART_CLK_M__L7_N0));
   INVX6M UART_CLK_M__L8_I1 (.Y(UART_CLK_M__L8_N1), 
	.A(UART_CLK_M__L7_N0));
   INVX6M UART_CLK_M__L8_I0 (.Y(UART_CLK_M__L8_N0), 
	.A(UART_CLK_M__L7_N0));
   CLKINVX32M UART_CLK_M__L7_I0 (.Y(UART_CLK_M__L7_N0), 
	.A(UART_CLK_M__L6_N0));
   CLKINVX40M UART_CLK_M__L6_I0 (.Y(UART_CLK_M__L6_N0), 
	.A(UART_CLK_M__L5_N0));
   CLKBUFX40M UART_CLK_M__L5_I0 (.Y(UART_CLK_M__L5_N0), 
	.A(UART_CLK_M__L4_N0));
   CLKBUFX40M UART_CLK_M__L4_I0 (.Y(UART_CLK_M__L4_N0), 
	.A(UART_CLK_M__L3_N0));
   CLKBUFX40M UART_CLK_M__L3_I0 (.Y(UART_CLK_M__L3_N0), 
	.A(UART_CLK_M__L2_N2));
   CLKBUFX40M UART_CLK_M__L2_I2 (.Y(UART_CLK_M__L2_N2), 
	.A(UART_CLK_M__L1_N0));
   INVX6M UART_CLK_M__L2_I1 (.Y(UART_CLK_M__L2_N1), 
	.A(UART_CLK_M__L1_N0));
   INVX6M UART_CLK_M__L2_I0 (.Y(UART_CLK_M__L2_N0), 
	.A(UART_CLK_M__L1_N0));
   CLKINVX24M UART_CLK_M__L1_I0 (.Y(UART_CLK_M__L1_N0), 
	.A(UART_CLK_M));
   CLKBUFX40M RX_CLK_M__L1_I0 (.Y(RX_CLK_M__L1_N0), 
	.A(RX_CLK_M));
   CLKBUFX40M TX_CLK_M__L1_I0 (.Y(TX_CLK_M__L1_N0), 
	.A(TX_CLK_M));
   BUFX4M FE_OFC24_SE (.Y(FE_OFN24_SE), 
	.A(FE_OFN17_SE));
   BUFX4M FE_OFC22_SE (.Y(FE_OFN22_SE), 
	.A(FE_OFN18_SE));
   CLKBUFX6M FE_OFC21_SE (.Y(FE_OFN21_SE), 
	.A(SE));
   BUFX4M FE_OFC20_SE (.Y(FE_OFN20_SE), 
	.A(SE));
   BUFX4M FE_OFC19_SE (.Y(FE_OFN19_SE), 
	.A(SE));
   BUFX4M FE_OFC18_SE (.Y(FE_OFN18_SE), 
	.A(SE));
   CLKBUFX6M FE_OFC17_SE (.Y(FE_OFN17_SE), 
	.A(SE));
   BUFX8M FE_OFC15_RST_D2_M (.Y(FE_OFN15_RST_D2_M), 
	.A(FE_OFN14_RST_D2_M));
   BUFX8M FE_OFC14_RST_D2_M (.Y(FE_OFN14_RST_D2_M), 
	.A(RST_D2_M));
   BUFX8M FE_OFC12_RST_D1_M (.Y(FE_OFN12_RST_D1_M), 
	.A(FE_OFN10_RST_D1_M));
   BUFX6M FE_OFC11_RST_D1_M (.Y(FE_OFN11_RST_D1_M), 
	.A(FE_OFN10_RST_D1_M));
   BUFX5M FE_OFC10_RST_D1_M (.Y(FE_OFN10_RST_D1_M), 
	.A(RST_D1_M));
   BUFX6M FE_OFC8_RST_D1_M (.Y(FE_OFN8_RST_D1_M), 
	.A(RST_D1_M));
   BUFX2M U4 (.Y(n1), 
	.A(Addr[0]));
   BUFX4M U5 (.Y(n2), 
	.A(Addr[1]));
   mux2X1_0 U0_mux2X1 (.IN_0(REF_CLK__L2_N0), 
	.IN_1(scan_clk__L3_N0), 
	.SEL(test_mode), 
	.OUT(REF_CLK_M));
   mux2X1_6 U1_mux2X1 (.IN_0(UART_CLK__L2_N0), 
	.IN_1(scan_clk__L2_N0), 
	.SEL(test_mode), 
	.OUT(UART_CLK_M));
   mux2X1_5 U2_mux2X1 (.IN_0(RST), 
	.IN_1(scan_rst), 
	.SEL(test_mode), 
	.OUT(RST_M));
   mux2X1_4 U3_mux2X1 (.IN_0(RX_CLK), 
	.IN_1(scan_clk__L5_N0), 
	.SEL(test_mode), 
	.OUT(RX_CLK_M));
   mux2X1_3 U4_mux2X1 (.IN_0(TX_CLK), 
	.IN_1(scan_clk__L5_N0), 
	.SEL(test_mode), 
	.OUT(TX_CLK_M));
   mux2X1_2 U5_mux2X1 (.IN_0(RST_D1), 
	.IN_1(scan_rst), 
	.SEL(test_mode), 
	.OUT(RST_D1_M));
   mux2X1_1 U6_mux2X1 (.IN_0(RST_D2), 
	.IN_1(scan_rst), 
	.SEL(test_mode), 
	.OUT(RST_D2_M));
   CLK_GATE CLK_GATE_dut (.E(Gate_En), 
	.CK(REF_CLK_M__L2_N0), 
	.test_en(test_mode), 
	.ECK(ALU_CLK));
   ClkDiv___test_1 CLK_DIV_TX_dut (.i_ref_clk(UART_CLK_M__L2_N0), 
	.i_rst_n(FE_OFN14_RST_D2_M), 
	.i_div_ratio({ 1'b0,
		1'b0,
		1'b1,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.o_div_clk(TX_CLK), 
	.test_si(n20), 
	.test_so(n19), 
	.test_se(SE), 
	.FE_OFN15_RST_D2_M(FE_OFN15_RST_D2_M), 
	.FE_OFN17_SE(FE_OFN17_SE), 
	.FE_OFN20_SE(FE_OFN20_SE), 
	.UART_CLK_M__L8_N0(UART_CLK_M__L8_N0), 
	.UART_CLK_M__L8_N2(UART_CLK_M__L8_N2), 
	.UART_CLK_M__L8_N3(UART_CLK_M__L8_N3));
   ClkDiv___test_0 CLK_DIV_RX_dut (.i_ref_clk(UART_CLK_M__L2_N1), 
	.i_rst_n(FE_OFN14_RST_D2_M), 
	.i_div_ratio({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b1,
		1'b0 }), 
	.o_div_clk(RX_CLK), 
	.test_si(n21), 
	.test_so(n20), 
	.test_se(FE_OFN17_SE), 
	.FE_OFN15_RST_D2_M(FE_OFN15_RST_D2_M), 
	.FE_OFN20_SE(FE_OFN20_SE), 
	.FE_OFN24_SE(FE_OFN24_SE), 
	.UART_CLK_M__L8_N0(UART_CLK_M__L8_N0), 
	.UART_CLK_M__L8_N1(UART_CLK_M__L8_N1), 
	.UART_CLK_M__L8_N2(UART_CLK_M__L8_N2));
   Rst_Sync_NUM_STAGES2_ACTIVE_TYPLOW_test_0 Rst_Sync_D1_dut (.RST(RST_M), 
	.CLK(REF_CLK_M__L5_N5), 
	.SYNC_RST(RST_D1), 
	.test_si(n13), 
	.test_so(n12), 
	.test_se(FE_OFN22_SE));
   Rst_Sync_NUM_STAGES2_ACTIVE_TYPLOW_test_1 Rst_Sync_D2_dut (.RST(RST_M), 
	.CLK(UART_CLK_M__L8_N3), 
	.SYNC_RST(RST_D2), 
	.test_si(n12), 
	.test_so(n11), 
	.test_se(SE), 
	.FE_OFN22_SE(FE_OFN22_SE));
   Data_Sync_NUM_STAGES2_BUS_WIDTH8_test_1 Data_Sync_dut (.CLK(REF_CLK_M__L5_N0), 
	.RST_n(FE_OFN10_RST_D1_M), 
	.bus_enable(in_Data_Sys_en), 
	.UNSYNC_bus({ in_Data_Sys[7],
		in_Data_Sys[6],
		in_Data_Sys[5],
		in_Data_Sys[4],
		in_Data_Sys[3],
		in_Data_Sys[2],
		in_Data_Sys[1],
		in_Data_Sys[0] }), 
	.enable_pulse(enable_pulse), 
	.SYNC_bus({ SYNC_bus[7],
		SYNC_bus[6],
		SYNC_bus[5],
		SYNC_bus[4],
		SYNC_bus[3],
		SYNC_bus[2],
		SYNC_bus[1],
		SYNC_bus[0] }), 
	.test_si2(test_si4), 
	.test_si1(n19), 
	.test_so2(n16), 
	.test_so1(test_so3), 
	.test_se(SE), 
	.FE_OFN8_RST_D1_M(FE_OFN8_RST_D1_M), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.REF_CLK_M__L5_N1(REF_CLK_M__L5_N1));
   SYS_CTRL_test_1 SYS_CTRL_dut (.CLK(REF_CLK_M__L5_N0), 
	.RST(FE_OFN10_RST_D1_M), 
	.Data_sync({ SYNC_bus[7],
		SYNC_bus[6],
		SYNC_bus[5],
		SYNC_bus[4],
		SYNC_bus[3],
		SYNC_bus[2],
		SYNC_bus[1],
		SYNC_bus[0] }), 
	.enable_pulse(enable_pulse), 
	.FIFO_FULL(F_Full), 
	.Rd_DATA({ RdData[7],
		RdData[6],
		RdData[5],
		RdData[4],
		RdData[3],
		RdData[2],
		RdData[1],
		RdData[0] }), 
	.Rd_Valid(Rd_Valid), 
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }), 
	.OUT_VALID(OUT_VALID), 
	.WR_DATA({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }), 
	.WR_INC(WR_INC), 
	.FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }), 
	.EN(Enable), 
	.Gate_En(Gate_En), 
	.Wr_D({ Wr_D[7],
		Wr_D[6],
		Wr_D[5],
		Wr_D[4],
		Wr_D[3],
		Wr_D[2],
		Wr_D[1],
		Wr_D[0] }), 
	.Addr({ SYNOPSYS_UNCONNECTED__0,
		SYNOPSYS_UNCONNECTED__1,
		SYNOPSYS_UNCONNECTED__2,
		SYNOPSYS_UNCONNECTED__3,
		Addr[3],
		Addr[2],
		Addr[1],
		Addr[0] }), 
	.RdEn(RdEn), 
	.WrEn(WrEn), 
	.test_si(n11), 
	.test_so(n10), 
	.test_se(SE), 
	.FE_OFN11_RST_D1_M(FE_OFN11_RST_D1_M), 
	.FE_OFN12_RST_D1_M(FE_OFN12_RST_D1_M), 
	.FE_OFN8_RST_D1_M(FE_OFN8_RST_D1_M), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.FE_OFN19_SE(FE_OFN19_SE), 
	.REF_CLK_M__L5_N1(REF_CLK_M__L5_N1), 
	.REF_CLK_M__L5_N2(REF_CLK_M__L5_N2));
   Register_File_10_0_1_test_1 Reg_file_dut (.CLK(REF_CLK_M__L5_N1), 
	.RST_n(RST_D1_M), 
	.RdEn(RdEn), 
	.WrEn(WrEn), 
	.Address({ Addr[3],
		Addr[2],
		n2,
		n1 }), 
	.WrData({ Wr_D[7],
		Wr_D[6],
		Wr_D[5],
		Wr_D[4],
		Wr_D[3],
		Wr_D[2],
		Wr_D[1],
		Wr_D[0] }), 
	.RdData({ RdData[7],
		RdData[6],
		RdData[5],
		RdData[4],
		RdData[3],
		RdData[2],
		RdData[1],
		RdData[0] }), 
	.RdData_Valid(Rd_Valid), 
	.REG0({ REG0[7],
		REG0[6],
		REG0[5],
		REG0[4],
		REG0[3],
		REG0[2],
		REG0[1],
		REG0[0] }), 
	.REG1({ REG1[7],
		REG1[6],
		REG1[5],
		REG1[4],
		REG1[3],
		REG1[2],
		REG1[1],
		REG1[0] }), 
	.REG3 (), 
	.test_si2(test_si5), 
	.test_si1(n16), 
	.test_so2(n13), 
	.test_so1(test_so4), 
	.test_se(SE), 
	.FE_OFN10_RST_D1_M(FE_OFN10_RST_D1_M), 
	.FE_OFN11_RST_D1_M(FE_OFN11_RST_D1_M), 
	.FE_OFN8_RST_D1_M(FE_OFN8_RST_D1_M), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.FE_OFN19_SE(FE_OFN19_SE), 
	.FE_OFN22_SE(FE_OFN22_SE), 
	.REF_CLK_M__L5_N2(REF_CLK_M__L5_N2), 
	.REF_CLK_M__L5_N5(REF_CLK_M__L5_N5), 
	.REF_CLK_M__L5_N6(REF_CLK_M__L5_N6));
   ALU_00000008_00000004_test_1 ALU_dut (.CLK(ALU_CLK__L1_N0), 
	.RST_n(FE_OFN11_RST_D1_M), 
	.A({ REG0[7],
		REG0[6],
		REG0[5],
		REG0[4],
		REG0[3],
		REG0[2],
		REG0[1],
		REG0[0] }), 
	.B({ REG1[7],
		REG1[6],
		REG1[5],
		REG1[4],
		REG1[3],
		REG1[2],
		REG1[1],
		REG1[0] }), 
	.ALU_FUN({ ALU_FUN[3],
		ALU_FUN[2],
		ALU_FUN[1],
		ALU_FUN[0] }), 
	.Enable(Enable), 
	.ALU_OUT({ ALU_OUT[15],
		ALU_OUT[14],
		ALU_OUT[13],
		ALU_OUT[12],
		ALU_OUT[11],
		ALU_OUT[10],
		ALU_OUT[9],
		ALU_OUT[8],
		ALU_OUT[7],
		ALU_OUT[6],
		ALU_OUT[5],
		ALU_OUT[4],
		ALU_OUT[3],
		ALU_OUT[2],
		ALU_OUT[1],
		ALU_OUT[0] }), 
	.OUT_VALID(OUT_VALID), 
	.test_si(SI), 
	.test_se(FE_OFN19_SE), 
	.FE_OFN12_RST_D1_M(FE_OFN12_RST_D1_M), 
	.FE_OFN21_SE(FE_OFN21_SE));
   UART_TX_test_1 UART_TX_dut (.CLK(TX_CLK_M__L1_N0), 
	.RST_n(FE_OFN15_RST_D2_M), 
	.P_DATA({ in_DATA_tx[7],
		in_DATA_tx[6],
		in_DATA_tx[5],
		in_DATA_tx[4],
		in_DATA_tx[3],
		in_DATA_tx[2],
		in_DATA_tx[1],
		in_DATA_tx[0] }), 
	.PAR_EN(1'b1), 
	.PAR_TYP(1'b0), 
	.DATA_VALID(F_Empty), 
	.TX_OUT(TX_OUT), 
	.Busy(busy), 
	.test_si(n9), 
	.test_so(n8), 
	.test_se(FE_OFN24_SE));
   UART_RX_10_test_1 UART_RX_dut (.CLK(RX_CLK_M__L1_N0), 
	.RST_n(RST_D2_M), 
	.PAR_TYP(1'b0), 
	.PAR_EN(1'b1), 
	.Prescale({ 1'b0,
		1'b1,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.RX_IN(RX_IN), 
	.P_DATA({ in_Data_Sys[7],
		in_Data_Sys[6],
		in_Data_Sys[5],
		in_Data_Sys[4],
		in_Data_Sys[3],
		in_Data_Sys[2],
		in_Data_Sys[1],
		in_Data_Sys[0] }), 
	.DATA_Valid(in_Data_Sys_en), 
	.test_si(n10), 
	.test_so(n9), 
	.test_se(SE), 
	.FE_OFN14_RST_D2_M(FE_OFN14_RST_D2_M), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.FE_OFN22_SE(FE_OFN22_SE));
   ASYNC_FIFO_test_1 ASYNC_FIFO_dut (.W_CLK(REF_CLK_M__L5_N0), 
	.W_RST(RST_D1_M), 
	.W_INC(WR_INC), 
	.R_CLK(TX_CLK_M__L1_N0), 
	.R_RST(FE_OFN15_RST_D2_M), 
	.R_INC(R_INC), 
	.WR_DATA({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }), 
	.FULL(F_Full), 
	.EMPTY(F_Empty), 
	.RD_DATA({ in_DATA_tx[7],
		in_DATA_tx[6],
		in_DATA_tx[5],
		in_DATA_tx[4],
		in_DATA_tx[3],
		in_DATA_tx[2],
		in_DATA_tx[1],
		in_DATA_tx[0] }), 
	.test_si3(test_si3), 
	.test_si2(test_si2), 
	.test_si1(OUT_VALID), 
	.test_so3(n21), 
	.test_so2(test_so2), 
	.test_so1(SO), 
	.test_se(SE), 
	.FE_OFN10_RST_D1_M(FE_OFN10_RST_D1_M), 
	.FE_OFN11_RST_D1_M(FE_OFN11_RST_D1_M), 
	.FE_OFN12_RST_D1_M(FE_OFN12_RST_D1_M), 
	.FE_OFN17_SE(FE_OFN17_SE), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.FE_OFN21_SE(FE_OFN21_SE), 
	.FE_OFN24_SE(FE_OFN24_SE), 
	.REF_CLK_M__L5_N2(REF_CLK_M__L5_N2), 
	.REF_CLK_M__L5_N3(REF_CLK_M__L5_N3), 
	.REF_CLK_M__L5_N4(REF_CLK_M__L5_N4), 
	.REF_CLK_M__L5_N7(REF_CLK_M__L5_N7));
   PULSE_GENERATOR_test_1 pulse_gen_dut (.CLK(TX_CLK_M__L1_N0), 
	.RST_n(FE_OFN15_RST_D2_M), 
	.in(busy), 
	.out(R_INC), 
	.test_si(n8), 
	.test_se(FE_OFN24_SE));
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Thu Sep 21 15:14:42 2023
/////////////////////////////////////////////////////////////
module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   AO2B2X4M U1 (.Y(OUT), 
	.B1(IN_1), 
	.B0(SEL), 
	.A1N(SEL), 
	.A0(IN_0));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   AO2B2X2M U1 (.Y(OUT), 
	.B1(IN_1), 
	.B0(SEL), 
	.A1N(SEL), 
	.A0(IN_0));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   AO2B2X2M U1 (.Y(OUT), 
	.B1(IN_1), 
	.B0(SEL), 
	.A1N(SEL), 
	.A0(IN_0));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   AO2B2X2M U1 (.Y(OUT), 
	.B1(IN_1), 
	.B0(SEL), 
	.A1N(SEL), 
	.A0(IN_0));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   AO2B2X2M U1 (.Y(OUT), 
	.B1(IN_1), 
	.B0(SEL), 
	.A1N(SEL), 
	.A0(IN_0));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   AO2B2X4M U1 (.Y(OUT), 
	.B1(IN_1), 
	.B0(SEL), 
	.A1N(SEL), 
	.A0(IN_0));
endmodule

module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;

   AO2B2X2M U1 (.Y(OUT), 
	.B1(IN_1), 
	.B0(SEL), 
	.A1N(SEL), 
	.A0(IN_0));
endmodule

module CLK_GATE (
	E, 
	CK, 
	test_en, 
	ECK);
   input E;
   input CK;
   input test_en;
   output ECK;

   // Internal wires
   wire _0_net_;

   TLATNCAX3M ICG_DUT (.ECK(ECK), 
	.E(_0_net_), 
	.CK(CK));
   OR2X2M U1 (.Y(_0_net_), 
	.B(test_en), 
	.A(E));
endmodule

module ClkDiv___0_DW01_inc_0 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___0_DW01_inc_1 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___0_DW01_inc_2 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___0_DW01_inc_3 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN15_RST_D2_M, 
	FE_OFN17_SE, 
	FE_OFN20_SE, 
	UART_CLK_M__L8_N0, 
	UART_CLK_M__L8_N2, 
	UART_CLK_M__L8_N3);
   input i_ref_clk;
   input i_rst_n;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN15_RST_D2_M;
   input FE_OFN17_SE;
   input FE_OFN20_SE;
   input UART_CLK_M__L8_N0;
   input UART_CLK_M__L8_N2;
   input UART_CLK_M__L8_N3;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire even_ratio_31;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N67;
   wire N162;
   wire n64;
   wire n65;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire \add_43/carry[7] ;
   wire \add_43/carry[6] ;
   wire \add_43/carry[5] ;
   wire \add_43/carry[4] ;
   wire \add_43/carry[3] ;
   wire \add_43/carry[2] ;
   wire n2;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n62;
   wire n63;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire [6:0] even_ratio;
   wire [31:0] half_low;
   wire [9:0] Counter_1;
   wire [9:0] Counter_2;
   wire [9:0] Counter_3;
   wire [9:0] Counter_4;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   SDFFRQX2M \current_state_reg[1]  (.SI(current_state[0]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(current_state[1]), 
	.D(next_state[1]), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \current_state_reg[0]  (.SI(Counter_4[9]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_4_reg[4]  (.SI(Counter_4[3]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[4]), 
	.D(n108), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_4_reg[6]  (.SI(Counter_4[5]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_4[6]), 
	.D(n106), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_3_reg[6]  (.SI(Counter_3[5]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_3[6]), 
	.D(n115), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_3_reg[4]  (.SI(Counter_3[3]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[4]), 
	.D(n117), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_1_reg[9]  (.SI(Counter_1[8]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[9]), 
	.D(n123), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[9]  (.SI(Counter_4[8]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_4[9]), 
	.D(n103), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_3_reg[9]  (.SI(Counter_3[8]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_3[9]), 
	.D(n122), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \current_state_reg[2]  (.SI(current_state[1]), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(current_state[2]), 
	.D(n186), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[9]  (.SI(Counter_2[8]), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[9]), 
	.D(n84), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_4_reg[0]  (.SI(Counter_3[9]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_4[0]), 
	.D(n112), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_3_reg[0]  (.SI(Counter_2[9]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[0]), 
	.D(n121), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_1_reg[0]  (.SI(test_si), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[0]), 
	.D(n102), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[0]  (.SI(Counter_1[9]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_2[0]), 
	.D(n93), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_1_reg[8]  (.SI(Counter_1[7]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[8]), 
	.D(n94), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[8]  (.SI(Counter_4[7]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_4[8]), 
	.D(n104), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_3_reg[8]  (.SI(Counter_3[7]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_3[8]), 
	.D(n113), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_4_reg[1]  (.SI(Counter_4[0]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_4[1]), 
	.D(n111), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_4_reg[2]  (.SI(Counter_4[1]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_4[2]), 
	.D(n110), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_4_reg[3]  (.SI(Counter_4[2]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[3]), 
	.D(n109), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_4_reg[5]  (.SI(Counter_4[4]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[5]), 
	.D(n107), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_3_reg[5]  (.SI(Counter_3[4]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[5]), 
	.D(n116), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_3_reg[3]  (.SI(Counter_3[2]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[3]), 
	.D(n118), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_3_reg[2]  (.SI(Counter_3[1]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[2]), 
	.D(n119), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_3_reg[1]  (.SI(Counter_3[0]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[1]), 
	.D(n120), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_4_reg[7]  (.SI(Counter_4[6]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_4[7]), 
	.D(n105), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_3_reg[7]  (.SI(Counter_3[6]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_3[7]), 
	.D(n114), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_1_reg[6]  (.SI(Counter_1[5]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[6]), 
	.D(n96), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_1_reg[4]  (.SI(Counter_1[3]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[4]), 
	.D(n98), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_1_reg[5]  (.SI(Counter_1[4]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[5]), 
	.D(n97), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_1_reg[3]  (.SI(Counter_1[2]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[3]), 
	.D(n99), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_1_reg[2]  (.SI(Counter_1[1]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[2]), 
	.D(n100), 
	.CK(UART_CLK_M__L8_N3));
   SDFFRQX2M \Counter_1_reg[1]  (.SI(Counter_1[0]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[1]), 
	.D(n101), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_2_reg[2]  (.SI(Counter_2[1]), 
	.SE(FE_OFN20_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[2]), 
	.D(n91), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[3]  (.SI(Counter_2[2]), 
	.SE(FE_OFN20_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[3]), 
	.D(n90), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[4]  (.SI(Counter_2[3]), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[4]), 
	.D(n89), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[5]  (.SI(Counter_2[4]), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[5]), 
	.D(n88), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[6]  (.SI(Counter_2[5]), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[6]), 
	.D(n87), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[7]  (.SI(Counter_2[6]), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[7]), 
	.D(n86), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[8]  (.SI(Counter_2[7]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_2[8]), 
	.D(n85), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_1_reg[7]  (.SI(Counter_1[6]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_1[7]), 
	.D(n95), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_2_reg[1]  (.SI(Counter_2[0]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_2[1]), 
	.D(n92), 
	.CK(UART_CLK_M__L8_N2));
   AOI31X2M U52 (.Y(n64), 
	.B0(n65), 
	.A2(n187), 
	.A1(n188), 
	.A0(i_ref_clk));
   NAND2X2M U12 (.Y(n142), 
	.B(n131), 
	.A(n83));
   NOR2X2M U51 (.Y(n2), 
	.B(n146), 
	.A(n143));
   NOR2X2M U53 (.Y(n148), 
	.B(n146), 
	.A(n143));
   INVX2M U54 (.Y(n146), 
	.A(n141));
   INVX2M U55 (.Y(n152), 
	.A(n83));
   INVX2M U56 (.Y(n150), 
	.A(n131));
   INVX2M U57 (.Y(n80), 
	.A(n66));
   INVX2M U62 (.Y(n143), 
	.A(n130));
   NAND2BX2M U63 (.Y(n66), 
	.B(even_ratio_31), 
	.AN(\add_43/carry[7] ));
   ADDHX1M U64 (.S(half_low[5]), 
	.CO(\add_43/carry[6] ), 
	.B(\add_43/carry[5] ), 
	.A(even_ratio[5]));
   ADDHX1M U65 (.S(half_low[2]), 
	.CO(\add_43/carry[3] ), 
	.B(\add_43/carry[2] ), 
	.A(even_ratio[2]));
   ADDHX1M U66 (.S(half_low[3]), 
	.CO(\add_43/carry[4] ), 
	.B(\add_43/carry[3] ), 
	.A(even_ratio[3]));
   ADDHX1M U67 (.S(half_low[1]), 
	.CO(\add_43/carry[2] ), 
	.B(even_ratio[0]), 
	.A(even_ratio[1]));
   ADDHX1M U68 (.S(half_low[4]), 
	.CO(\add_43/carry[5] ), 
	.B(\add_43/carry[4] ), 
	.A(even_ratio[4]));
   ADDHX1M U69 (.S(half_low[6]), 
	.CO(\add_43/carry[7] ), 
	.B(\add_43/carry[6] ), 
	.A(even_ratio[6]));
   OR2X2M U73 (.Y(n10), 
	.B(LTIE_LTIELO_NET), 
	.A(LTIE_LTIELO_NET));
   CLKINVX1M U74 (.Y(even_ratio[0]), 
	.A(LTIE_LTIELO_NET));
   OAI2BB1X1M U75 (.Y(even_ratio[1]), 
	.B0(n10), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(LTIE_LTIELO_NET));
   OR2X1M U76 (.Y(n11), 
	.B(LTIE_LTIELO_NET), 
	.A(n10));
   OAI2BB1X1M U77 (.Y(even_ratio[2]), 
	.B0(n11), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(n10));
   OR2X1M U78 (.Y(n12), 
	.B(LTIE_LTIELO_NET), 
	.A(n11));
   OAI2BB1X1M U79 (.Y(even_ratio[3]), 
	.B0(n12), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(n11));
   OR2X1M U80 (.Y(n13), 
	.B(HTIE_LTIEHI_NET), 
	.A(n12));
   OAI2BB1X1M U81 (.Y(even_ratio[4]), 
	.B0(n13), 
	.A1N(HTIE_LTIEHI_NET), 
	.A0N(n12));
   XNOR2X1M U82 (.Y(even_ratio[5]), 
	.B(n13), 
	.A(LTIE_LTIELO_NET));
   NOR3X1M U83 (.Y(even_ratio_31), 
	.C(n13), 
	.B(LTIE_LTIELO_NET), 
	.A(LTIE_LTIELO_NET));
   OAI21X1M U84 (.Y(n14), 
	.B0(LTIE_LTIELO_NET), 
	.A1(n13), 
	.A0(LTIE_LTIELO_NET));
   NAND2BX1M U85 (.Y(even_ratio[6]), 
	.B(n14), 
	.AN(even_ratio_31));
   CLKXOR2X2M U86 (.Y(half_low[7]), 
	.B(even_ratio_31), 
	.A(\add_43/carry[7] ));
   NOR2BX1M U88 (.Y(n62), 
	.B(Counter_2[0]), 
	.AN(LTIE_LTIELO_NET));
   OAI2B2X1M U89 (.Y(n68), 
	.B1(n62), 
	.B0(half_low[1]), 
	.A1N(Counter_2[1]), 
	.A0(n62));
   NOR2BX1M U90 (.Y(n63), 
	.B(LTIE_LTIELO_NET), 
	.AN(Counter_2[0]));
   OAI2B2X1M U91 (.Y(n67), 
	.B1(n63), 
	.B0(Counter_2[1]), 
	.A1N(half_low[1]), 
	.A0(n63));
   XNOR2X1M U93 (.Y(n72), 
	.B(Counter_2[5]), 
	.A(half_low[5]));
   XNOR2X1M U94 (.Y(n71), 
	.B(Counter_2[4]), 
	.A(half_low[4]));
   XNOR2X1M U95 (.Y(n70), 
	.B(Counter_2[3]), 
	.A(half_low[3]));
   XNOR2X1M U96 (.Y(n69), 
	.B(Counter_2[2]), 
	.A(half_low[2]));
   NAND4X1M U97 (.Y(n78), 
	.D(n69), 
	.C(n70), 
	.B(n71), 
	.A(n72));
   XNOR2X1M U98 (.Y(n76), 
	.B(Counter_2[9]), 
	.A(n80));
   XNOR2X1M U99 (.Y(n75), 
	.B(Counter_2[8]), 
	.A(n80));
   XNOR2X1M U100 (.Y(n74), 
	.B(Counter_2[7]), 
	.A(half_low[7]));
   XNOR2X1M U101 (.Y(n73), 
	.B(Counter_2[6]), 
	.A(half_low[6]));
   NAND4X1M U102 (.Y(n77), 
	.D(n73), 
	.C(n74), 
	.B(n75), 
	.A(n76));
   NOR4X1M U103 (.Y(N162), 
	.D(n77), 
	.C(n78), 
	.B(n79), 
	.A(n80));
   CLKINVX1M U104 (.Y(o_div_clk), 
	.A(n64));
   OAI211X1M U105 (.Y(next_state[1]), 
	.C0(n124), 
	.B0(n83), 
	.A1(n82), 
	.A0(n81));
   AOI2B1X1M U106 (.Y(n124), 
	.B0(n127), 
	.A1N(n125), 
	.A0(n126));
   AOI21X1M U107 (.Y(n81), 
	.B0(n129), 
	.A1(n128), 
	.A0(n65));
   NAND4X1M U108 (.Y(next_state[0]), 
	.D(n133), 
	.C(n132), 
	.B(n131), 
	.A(n130));
   AOI221XLM U109 (.Y(n133), 
	.C0(n127), 
	.B1(n82), 
	.B0(n134), 
	.A1(n187), 
	.A0(n129));
   OAI2BB1X1M U110 (.Y(n127), 
	.B0(n135), 
	.A1N(N162), 
	.A0N(n134));
   OAI21X1M U111 (.Y(n135), 
	.B0(LTIE_LTIELO_NET), 
	.A1(n136), 
	.A0(n126));
   NOR3X1M U112 (.Y(n129), 
	.C(current_state[0]), 
	.B(current_state[2]), 
	.A(n137));
   NOR4BX1M U113 (.Y(n137), 
	.D(LTIE_LTIELO_NET), 
	.C(LTIE_LTIELO_NET), 
	.B(LTIE_LTIELO_NET), 
	.AN(n138));
   NOR4X1M U114 (.Y(n138), 
	.D(LTIE_LTIELO_NET), 
	.C(HTIE_LTIEHI_NET), 
	.B(LTIE_LTIELO_NET), 
	.A(LTIE_LTIELO_NET));
   NAND2BX1M U115 (.Y(n132), 
	.B(n136), 
	.AN(n139));
   OAI32X1M U116 (.Y(n186), 
	.B1(n141), 
	.B0(n82), 
	.A2(n140), 
	.A1(n187), 
	.A0(n128));
   CLKINVX1M U117 (.Y(n82), 
	.A(LTIE_LTIELO_NET));
   AO22X1M U118 (.Y(n99), 
	.B1(n143), 
	.B0(N28), 
	.A1(Counter_1[3]), 
	.A0(n142));
   AO22X1M U119 (.Y(n98), 
	.B1(n143), 
	.B0(N29), 
	.A1(Counter_1[4]), 
	.A0(n142));
   AO22X1M U120 (.Y(n97), 
	.B1(n143), 
	.B0(N30), 
	.A1(Counter_1[5]), 
	.A0(n142));
   AO22X1M U121 (.Y(n96), 
	.B1(n143), 
	.B0(N31), 
	.A1(Counter_1[6]), 
	.A0(n142));
   AO22X1M U122 (.Y(n95), 
	.B1(n143), 
	.B0(N32), 
	.A1(Counter_1[7]), 
	.A0(n142));
   OAI2BB2X1M U123 (.Y(n94), 
	.B1(n145), 
	.B0(n144), 
	.A1N(n143), 
	.A0N(N33));
   AO22X1M U124 (.Y(n93), 
	.B1(n146), 
	.B0(N36), 
	.A1(n142), 
	.A0(Counter_2[0]));
   AO22X1M U125 (.Y(n92), 
	.B1(n146), 
	.B0(N37), 
	.A1(n142), 
	.A0(Counter_2[1]));
   AO22X1M U126 (.Y(n91), 
	.B1(n146), 
	.B0(N38), 
	.A1(n142), 
	.A0(Counter_2[2]));
   AO22X1M U127 (.Y(n90), 
	.B1(n146), 
	.B0(N39), 
	.A1(n142), 
	.A0(Counter_2[3]));
   AO22X1M U128 (.Y(n89), 
	.B1(n146), 
	.B0(N40), 
	.A1(n142), 
	.A0(Counter_2[4]));
   AO22X1M U129 (.Y(n88), 
	.B1(n146), 
	.B0(N41), 
	.A1(n142), 
	.A0(Counter_2[5]));
   AO22X1M U130 (.Y(n87), 
	.B1(n146), 
	.B0(N42), 
	.A1(n142), 
	.A0(Counter_2[6]));
   AO22X1M U131 (.Y(n86), 
	.B1(n146), 
	.B0(N43), 
	.A1(n142), 
	.A0(Counter_2[7]));
   AO22X1M U132 (.Y(n85), 
	.B1(n146), 
	.B0(N44), 
	.A1(n142), 
	.A0(Counter_2[8]));
   AO22X1M U133 (.Y(n84), 
	.B1(n146), 
	.B0(N45), 
	.A1(n142), 
	.A0(Counter_2[9]));
   OAI2BB2X1M U134 (.Y(n123), 
	.B1(n147), 
	.B0(n144), 
	.A1N(n143), 
	.A0N(N34));
   CLKINVX1M U135 (.Y(n144), 
	.A(n142));
   OAI2BB2X1M U136 (.Y(n122), 
	.B1(n149), 
	.B0(n148), 
	.A1N(n150), 
	.A0N(N56));
   AO2B2X1M U137 (.Y(n121), 
	.B1(n150), 
	.B0(N47), 
	.A1N(n148), 
	.A0(Counter_3[0]));
   AO2B2X1M U138 (.Y(n120), 
	.B1(n150), 
	.B0(N48), 
	.A1N(n2), 
	.A0(Counter_3[1]));
   AO2B2X1M U139 (.Y(n119), 
	.B1(n150), 
	.B0(N49), 
	.A1N(n148), 
	.A0(Counter_3[2]));
   AO2B2X1M U140 (.Y(n118), 
	.B1(n150), 
	.B0(N50), 
	.A1N(n2), 
	.A0(Counter_3[3]));
   AO2B2X1M U141 (.Y(n117), 
	.B1(n150), 
	.B0(N51), 
	.A1N(n148), 
	.A0(Counter_3[4]));
   AO2B2X1M U142 (.Y(n116), 
	.B1(n150), 
	.B0(N52), 
	.A1N(n2), 
	.A0(Counter_3[5]));
   AO2B2X1M U143 (.Y(n115), 
	.B1(n150), 
	.B0(N53), 
	.A1N(n148), 
	.A0(Counter_3[6]));
   AO2B2X1M U144 (.Y(n114), 
	.B1(n150), 
	.B0(N54), 
	.A1N(n2), 
	.A0(Counter_3[7]));
   OAI2BB2X1M U145 (.Y(n113), 
	.B1(n151), 
	.B0(n2), 
	.A1N(n150), 
	.A0N(N55));
   AO2B2X1M U146 (.Y(n112), 
	.B1(n152), 
	.B0(N58), 
	.A1N(n148), 
	.A0(Counter_4[0]));
   AO2B2X1M U147 (.Y(n111), 
	.B1(n152), 
	.B0(N59), 
	.A1N(n2), 
	.A0(Counter_4[1]));
   AO2B2X1M U148 (.Y(n110), 
	.B1(n152), 
	.B0(N60), 
	.A1N(n148), 
	.A0(Counter_4[2]));
   AO2B2X1M U149 (.Y(n109), 
	.B1(n152), 
	.B0(N61), 
	.A1N(n2), 
	.A0(Counter_4[3]));
   AO2B2X1M U150 (.Y(n108), 
	.B1(n152), 
	.B0(N62), 
	.A1N(n148), 
	.A0(Counter_4[4]));
   AO2B2X1M U151 (.Y(n107), 
	.B1(n152), 
	.B0(N63), 
	.A1N(n2), 
	.A0(Counter_4[5]));
   AO2B2X1M U152 (.Y(n106), 
	.B1(n152), 
	.B0(N64), 
	.A1N(n148), 
	.A0(Counter_4[6]));
   AO2B2X1M U153 (.Y(n105), 
	.B1(n152), 
	.B0(N65), 
	.A1N(n2), 
	.A0(Counter_4[7]));
   OAI2BB2X1M U154 (.Y(n104), 
	.B1(n153), 
	.B0(n148), 
	.A1N(n152), 
	.A0N(N66));
   OAI2BB2X1M U155 (.Y(n103), 
	.B1(n154), 
	.B0(n2), 
	.A1N(n152), 
	.A0N(N67));
   NAND2BX1M U156 (.Y(n141), 
	.B(n134), 
	.AN(N162));
   NOR3X1M U157 (.Y(n134), 
	.C(n188), 
	.B(current_state[1]), 
	.A(current_state[0]));
   AO22X1M U158 (.Y(n102), 
	.B1(n143), 
	.B0(N25), 
	.A1(Counter_1[0]), 
	.A0(n142));
   AO22X1M U159 (.Y(n101), 
	.B1(n143), 
	.B0(N26), 
	.A1(Counter_1[1]), 
	.A0(n142));
   AO22X1M U160 (.Y(n100), 
	.B1(n143), 
	.B0(N27), 
	.A1(Counter_1[2]), 
	.A0(n142));
   NAND3X1M U161 (.Y(n130), 
	.C(n65), 
	.B(current_state[1]), 
	.A(n128));
   CLKINVX1M U162 (.Y(n65), 
	.A(n140));
   NAND4X1M U163 (.Y(n128), 
	.D(n158), 
	.C(n157), 
	.B(n156), 
	.A(n155));
   NOR4X1M U164 (.Y(n158), 
	.D(n161), 
	.C(Counter_1[7]), 
	.B(n160), 
	.A(n159));
   CLKXOR2X2M U165 (.Y(n161), 
	.B(Counter_1[0]), 
	.A(even_ratio[0]));
   CLKXOR2X2M U166 (.Y(n160), 
	.B(Counter_1[5]), 
	.A(even_ratio[5]));
   NAND3X1M U167 (.Y(n159), 
	.C(n145), 
	.B(n162), 
	.A(n147));
   CLKINVX1M U168 (.Y(n145), 
	.A(Counter_1[8]));
   CLKINVX1M U169 (.Y(n147), 
	.A(Counter_1[9]));
   NOR3X1M U170 (.Y(n157), 
	.C(n165), 
	.B(n164), 
	.A(n163));
   CLKXOR2X2M U171 (.Y(n165), 
	.B(Counter_1[1]), 
	.A(even_ratio[1]));
   CLKXOR2X2M U172 (.Y(n164), 
	.B(Counter_1[3]), 
	.A(even_ratio[3]));
   CLKXOR2X2M U173 (.Y(n163), 
	.B(Counter_1[2]), 
	.A(even_ratio[2]));
   XNOR2X1M U174 (.Y(n156), 
	.B(even_ratio[4]), 
	.A(Counter_1[4]));
   XNOR2X1M U175 (.Y(n155), 
	.B(even_ratio[6]), 
	.A(Counter_1[6]));
   CLKNAND2X2M U176 (.Y(n131), 
	.B(n125), 
	.A(n126));
   NAND4X1M U177 (.Y(n125), 
	.D(n169), 
	.C(n168), 
	.B(n167), 
	.A(n166));
   NOR4X1M U178 (.Y(n169), 
	.D(n172), 
	.C(Counter_3[7]), 
	.B(n171), 
	.A(n170));
   CLKXOR2X2M U179 (.Y(n172), 
	.B(Counter_3[0]), 
	.A(even_ratio[0]));
   CLKXOR2X2M U180 (.Y(n171), 
	.B(Counter_3[5]), 
	.A(even_ratio[5]));
   NAND3X1M U181 (.Y(n170), 
	.C(n151), 
	.B(n162), 
	.A(n149));
   CLKINVX1M U182 (.Y(n151), 
	.A(Counter_3[8]));
   CLKINVX1M U183 (.Y(n149), 
	.A(Counter_3[9]));
   NOR3X1M U184 (.Y(n168), 
	.C(n175), 
	.B(n174), 
	.A(n173));
   CLKXOR2X2M U185 (.Y(n175), 
	.B(Counter_3[1]), 
	.A(even_ratio[1]));
   CLKXOR2X2M U186 (.Y(n174), 
	.B(Counter_3[3]), 
	.A(even_ratio[3]));
   CLKXOR2X2M U187 (.Y(n173), 
	.B(Counter_3[2]), 
	.A(even_ratio[2]));
   XNOR2X1M U188 (.Y(n167), 
	.B(even_ratio[4]), 
	.A(Counter_3[4]));
   XNOR2X1M U189 (.Y(n166), 
	.B(even_ratio[6]), 
	.A(Counter_3[6]));
   NOR2X1M U190 (.Y(n126), 
	.B(current_state[1]), 
	.A(n140));
   CLKNAND2X2M U191 (.Y(n140), 
	.B(n188), 
	.A(current_state[0]));
   CLKINVX1M U192 (.Y(n188), 
	.A(current_state[2]));
   CLKNAND2X2M U193 (.Y(n83), 
	.B(n139), 
	.A(n136));
   NAND4X1M U194 (.Y(n139), 
	.D(n179), 
	.C(n178), 
	.B(n177), 
	.A(n176));
   NOR4X1M U195 (.Y(n179), 
	.D(n182), 
	.C(Counter_4[7]), 
	.B(n181), 
	.A(n180));
   CLKXOR2X2M U196 (.Y(n182), 
	.B(Counter_4[0]), 
	.A(even_ratio[0]));
   CLKXOR2X2M U197 (.Y(n181), 
	.B(Counter_4[5]), 
	.A(even_ratio[5]));
   NAND3X1M U198 (.Y(n180), 
	.C(n153), 
	.B(n162), 
	.A(n154));
   CLKINVX1M U199 (.Y(n153), 
	.A(Counter_4[8]));
   CLKINVX1M U200 (.Y(n162), 
	.A(even_ratio_31));
   CLKINVX1M U201 (.Y(n154), 
	.A(Counter_4[9]));
   NOR3X1M U202 (.Y(n178), 
	.C(n185), 
	.B(n184), 
	.A(n183));
   CLKXOR2X2M U203 (.Y(n185), 
	.B(Counter_4[1]), 
	.A(even_ratio[1]));
   CLKXOR2X2M U204 (.Y(n184), 
	.B(Counter_4[3]), 
	.A(even_ratio[3]));
   CLKXOR2X2M U205 (.Y(n183), 
	.B(Counter_4[2]), 
	.A(even_ratio[2]));
   XNOR2X1M U206 (.Y(n177), 
	.B(even_ratio[4]), 
	.A(Counter_4[4]));
   XNOR2X1M U207 (.Y(n176), 
	.B(even_ratio[6]), 
	.A(Counter_4[6]));
   NOR3X1M U208 (.Y(n136), 
	.C(n187), 
	.B(current_state[2]), 
	.A(current_state[0]));
   CLKINVX1M U209 (.Y(n187), 
	.A(current_state[1]));
   ClkDiv___0_DW01_inc_0 add_72 (.A({ Counter_4[9],
		Counter_4[8],
		Counter_4[7],
		Counter_4[6],
		Counter_4[5],
		Counter_4[4],
		Counter_4[3],
		Counter_4[2],
		Counter_4[1],
		Counter_4[0] }), 
	.SUM({ N67,
		N66,
		N65,
		N64,
		N63,
		N62,
		N61,
		N60,
		N59,
		N58 }));
   ClkDiv___0_DW01_inc_1 add_67 (.A({ Counter_3[9],
		Counter_3[8],
		Counter_3[7],
		Counter_3[6],
		Counter_3[5],
		Counter_3[4],
		Counter_3[3],
		Counter_3[2],
		Counter_3[1],
		Counter_3[0] }), 
	.SUM({ N56,
		N55,
		N54,
		N53,
		N52,
		N51,
		N50,
		N49,
		N48,
		N47 }));
   ClkDiv___0_DW01_inc_2 add_62 (.A({ Counter_2[9],
		Counter_2[8],
		Counter_2[7],
		Counter_2[6],
		Counter_2[5],
		Counter_2[4],
		Counter_2[3],
		Counter_2[2],
		Counter_2[1],
		Counter_2[0] }), 
	.SUM({ N45,
		N44,
		N43,
		N42,
		N41,
		N40,
		N39,
		N38,
		N37,
		N36 }));
   ClkDiv___0_DW01_inc_3 add_57 (.A({ Counter_1[9],
		Counter_1[8],
		Counter_1[7],
		Counter_1[6],
		Counter_1[5],
		Counter_1[4],
		Counter_1[3],
		Counter_1[2],
		Counter_1[1],
		Counter_1[0] }), 
	.SUM({ N34,
		N33,
		N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26,
		N25 }));
   NAND3BX2M U3 (.Y(n79), 
	.C(n68), 
	.B(n67), 
	.AN(n80));
endmodule

module ClkDiv___1_DW01_inc_0 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___1_DW01_inc_1 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___1_DW01_inc_2 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___1_DW01_inc_3 (
	A, 
	SUM);
   input [9:0] A;
   output [9:0] SUM;

   // Internal wires
   wire [9:2] carry;

   ADDHX1M U1_1_8 (.S(SUM[8]), 
	.CO(carry[9]), 
	.B(carry[8]), 
	.A(A[8]));
   ADDHX1M U1_1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.B(carry[6]), 
	.A(A[6]));
   ADDHX1M U1_1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.B(carry[4]), 
	.A(A[4]));
   ADDHX1M U1_1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.B(carry[5]), 
	.A(A[5]));
   ADDHX1M U1_1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.B(carry[3]), 
	.A(A[3]));
   ADDHX1M U1_1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.B(carry[2]), 
	.A(A[2]));
   ADDHX1M U1_1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.B(A[0]), 
	.A(A[1]));
   ADDHX1M U1_1_7 (.S(SUM[7]), 
	.CO(carry[8]), 
	.B(carry[7]), 
	.A(A[7]));
   CLKXOR2X2M U1 (.Y(SUM[9]), 
	.B(A[9]), 
	.A(carry[9]));
   CLKINVX1M U2 (.Y(SUM[0]), 
	.A(A[0]));
endmodule

module ClkDiv___test_0 (
	i_ref_clk, 
	i_rst_n, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN15_RST_D2_M, 
	FE_OFN20_SE, 
	FE_OFN24_SE, 
	UART_CLK_M__L8_N0, 
	UART_CLK_M__L8_N1, 
	UART_CLK_M__L8_N2);
   input i_ref_clk;
   input i_rst_n;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN15_RST_D2_M;
   input FE_OFN20_SE;
   input FE_OFN24_SE;
   input UART_CLK_M__L8_N0;
   input UART_CLK_M__L8_N1;
   input UART_CLK_M__L8_N2;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire even_ratio_31;
   wire N25;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire N65;
   wire N66;
   wire N67;
   wire N162;
   wire \add_43/carry[7] ;
   wire \add_43/carry[6] ;
   wire \add_43/carry[5] ;
   wire \add_43/carry[4] ;
   wire \add_43/carry[3] ;
   wire \add_43/carry[2] ;
   wire n2;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n62;
   wire n63;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire [6:0] even_ratio;
   wire [31:0] half_low;
   wire [9:0] Counter_1;
   wire [9:0] Counter_2;
   wire [9:0] Counter_3;
   wire [9:0] Counter_4;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = current_state[2] ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   SDFFRQX2M \current_state_reg[1]  (.SI(current_state[0]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(current_state[1]), 
	.D(next_state[1]), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \current_state_reg[0]  (.SI(Counter_4[9]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_4_reg[4]  (.SI(Counter_4[3]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[4]), 
	.D(n204), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[6]  (.SI(Counter_4[5]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[6]), 
	.D(n206), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[6]  (.SI(Counter_3[5]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[6]), 
	.D(n197), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[4]  (.SI(Counter_3[3]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[4]), 
	.D(n195), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_1_reg[9]  (.SI(Counter_1[8]), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[9]), 
	.D(n189), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_4_reg[9]  (.SI(Counter_4[8]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_4[9]), 
	.D(n209), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_3_reg[9]  (.SI(Counter_3[8]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[9]), 
	.D(n190), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \current_state_reg[2]  (.SI(current_state[1]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(current_state[2]), 
	.D(n186), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[9]  (.SI(Counter_2[8]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_2[9]), 
	.D(n228), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_4_reg[0]  (.SI(Counter_3[9]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[0]), 
	.D(n200), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[0]  (.SI(Counter_2[9]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_3[0]), 
	.D(n191), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_1_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[0]), 
	.D(n210), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[0]  (.SI(Counter_1[9]), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[0]), 
	.D(n219), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_1_reg[8]  (.SI(Counter_1[7]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[8]), 
	.D(n218), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_4_reg[8]  (.SI(Counter_4[7]), 
	.SE(FE_OFN20_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_4[8]), 
	.D(n208), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[8]  (.SI(Counter_3[7]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[8]), 
	.D(n199), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[1]  (.SI(Counter_4[0]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[1]), 
	.D(n201), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[2]  (.SI(Counter_4[1]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[2]), 
	.D(n202), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[3]  (.SI(Counter_4[2]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[3]), 
	.D(n203), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[5]  (.SI(Counter_4[4]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[5]), 
	.D(n205), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[5]  (.SI(Counter_3[4]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[5]), 
	.D(n196), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[3]  (.SI(Counter_3[2]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[3]), 
	.D(n194), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[2]  (.SI(Counter_3[1]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_3[2]), 
	.D(n193), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_3_reg[1]  (.SI(Counter_3[0]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[1]), 
	.D(n192), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_4_reg[7]  (.SI(Counter_4[6]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_4[7]), 
	.D(n207), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_3_reg[7]  (.SI(Counter_3[6]), 
	.SE(FE_OFN20_SE), 
	.RN(i_rst_n), 
	.Q(Counter_3[7]), 
	.D(n198), 
	.CK(UART_CLK_M__L8_N2));
   SDFFRQX2M \Counter_1_reg[6]  (.SI(Counter_1[5]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[6]), 
	.D(n216), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_1_reg[4]  (.SI(Counter_1[3]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[4]), 
	.D(n214), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_1_reg[5]  (.SI(Counter_1[4]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[5]), 
	.D(n215), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_1_reg[3]  (.SI(Counter_1[2]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[3]), 
	.D(n213), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_1_reg[2]  (.SI(Counter_1[1]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[2]), 
	.D(n212), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_1_reg[1]  (.SI(Counter_1[0]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[1]), 
	.D(n211), 
	.CK(UART_CLK_M__L8_N0));
   SDFFRQX2M \Counter_2_reg[2]  (.SI(Counter_2[1]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[2]), 
	.D(n221), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_2_reg[3]  (.SI(Counter_2[2]), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[3]), 
	.D(n222), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_2_reg[4]  (.SI(Counter_2[3]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[4]), 
	.D(n223), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_2_reg[5]  (.SI(Counter_2[4]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[5]), 
	.D(n224), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_2_reg[6]  (.SI(Counter_2[5]), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[6]), 
	.D(n225), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_2_reg[7]  (.SI(Counter_2[6]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_2[7]), 
	.D(n226), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_2_reg[8]  (.SI(Counter_2[7]), 
	.SE(test_se), 
	.RN(i_rst_n), 
	.Q(Counter_2[8]), 
	.D(n227), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_1_reg[7]  (.SI(Counter_1[6]), 
	.SE(test_se), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_1[7]), 
	.D(n217), 
	.CK(UART_CLK_M__L8_N1));
   SDFFRQX2M \Counter_2_reg[1]  (.SI(Counter_2[0]), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN15_RST_D2_M), 
	.Q(Counter_2[1]), 
	.D(n220), 
	.CK(UART_CLK_M__L8_N1));
   AOI31X2M U52 (.Y(n230), 
	.B0(n229), 
	.A2(n187), 
	.A1(n188), 
	.A0(i_ref_clk));
   NAND2X2M U12 (.Y(n142), 
	.B(n131), 
	.A(n83));
   NOR2X2M U51 (.Y(n2), 
	.B(n146), 
	.A(n143));
   NOR2X2M U53 (.Y(n148), 
	.B(n146), 
	.A(n143));
   INVX2M U54 (.Y(n146), 
	.A(n141));
   INVX2M U55 (.Y(n152), 
	.A(n83));
   INVX2M U56 (.Y(n150), 
	.A(n131));
   INVX2M U57 (.Y(n80), 
	.A(n66));
   INVX2M U62 (.Y(n143), 
	.A(n130));
   NAND2BX2M U63 (.Y(n66), 
	.B(even_ratio_31), 
	.AN(\add_43/carry[7] ));
   ADDHX1M U64 (.S(half_low[5]), 
	.CO(\add_43/carry[6] ), 
	.B(\add_43/carry[5] ), 
	.A(even_ratio[5]));
   ADDHX1M U65 (.S(half_low[2]), 
	.CO(\add_43/carry[3] ), 
	.B(\add_43/carry[2] ), 
	.A(even_ratio[2]));
   ADDHX1M U66 (.S(half_low[3]), 
	.CO(\add_43/carry[4] ), 
	.B(\add_43/carry[3] ), 
	.A(even_ratio[3]));
   ADDHX1M U67 (.S(half_low[1]), 
	.CO(\add_43/carry[2] ), 
	.B(even_ratio[0]), 
	.A(even_ratio[1]));
   ADDHX1M U68 (.S(half_low[4]), 
	.CO(\add_43/carry[5] ), 
	.B(\add_43/carry[4] ), 
	.A(even_ratio[4]));
   ADDHX1M U69 (.S(half_low[6]), 
	.CO(\add_43/carry[7] ), 
	.B(\add_43/carry[6] ), 
	.A(even_ratio[6]));
   OR2X2M U73 (.Y(n10), 
	.B(HTIE_LTIEHI_NET), 
	.A(LTIE_LTIELO_NET));
   CLKINVX1M U74 (.Y(even_ratio[0]), 
	.A(HTIE_LTIEHI_NET));
   OAI2BB1X1M U75 (.Y(even_ratio[1]), 
	.B0(n10), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(HTIE_LTIEHI_NET));
   OR2X1M U76 (.Y(n11), 
	.B(LTIE_LTIELO_NET), 
	.A(n10));
   OAI2BB1X1M U77 (.Y(even_ratio[2]), 
	.B0(n11), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(n10));
   OR2X1M U78 (.Y(n12), 
	.B(LTIE_LTIELO_NET), 
	.A(n11));
   OAI2BB1X1M U79 (.Y(even_ratio[3]), 
	.B0(n12), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(n11));
   OR2X1M U80 (.Y(n13), 
	.B(LTIE_LTIELO_NET), 
	.A(n12));
   OAI2BB1X1M U81 (.Y(even_ratio[4]), 
	.B0(n13), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(n12));
   XNOR2X1M U82 (.Y(even_ratio[5]), 
	.B(n13), 
	.A(LTIE_LTIELO_NET));
   NOR3X1M U83 (.Y(even_ratio_31), 
	.C(n13), 
	.B(LTIE_LTIELO_NET), 
	.A(LTIE_LTIELO_NET));
   OAI21X1M U84 (.Y(n14), 
	.B0(LTIE_LTIELO_NET), 
	.A1(n13), 
	.A0(LTIE_LTIELO_NET));
   NAND2BX1M U85 (.Y(even_ratio[6]), 
	.B(n14), 
	.AN(even_ratio_31));
   CLKXOR2X2M U86 (.Y(half_low[7]), 
	.B(even_ratio_31), 
	.A(\add_43/carry[7] ));
   NOR2BX1M U88 (.Y(n62), 
	.B(Counter_2[0]), 
	.AN(HTIE_LTIEHI_NET));
   OAI2B2X1M U89 (.Y(n68), 
	.B1(n62), 
	.B0(half_low[1]), 
	.A1N(Counter_2[1]), 
	.A0(n62));
   NOR2BX1M U90 (.Y(n63), 
	.B(HTIE_LTIEHI_NET), 
	.AN(Counter_2[0]));
   OAI2B2X1M U91 (.Y(n67), 
	.B1(n63), 
	.B0(Counter_2[1]), 
	.A1N(half_low[1]), 
	.A0(n63));
   XNOR2X1M U93 (.Y(n72), 
	.B(Counter_2[5]), 
	.A(half_low[5]));
   XNOR2X1M U94 (.Y(n71), 
	.B(Counter_2[4]), 
	.A(half_low[4]));
   XNOR2X1M U95 (.Y(n70), 
	.B(Counter_2[3]), 
	.A(half_low[3]));
   XNOR2X1M U96 (.Y(n69), 
	.B(Counter_2[2]), 
	.A(half_low[2]));
   NAND4X1M U97 (.Y(n78), 
	.D(n69), 
	.C(n70), 
	.B(n71), 
	.A(n72));
   XNOR2X1M U98 (.Y(n76), 
	.B(Counter_2[9]), 
	.A(n80));
   XNOR2X1M U99 (.Y(n75), 
	.B(Counter_2[8]), 
	.A(n80));
   XNOR2X1M U100 (.Y(n74), 
	.B(Counter_2[7]), 
	.A(half_low[7]));
   XNOR2X1M U101 (.Y(n73), 
	.B(Counter_2[6]), 
	.A(half_low[6]));
   NAND4X1M U102 (.Y(n77), 
	.D(n73), 
	.C(n74), 
	.B(n75), 
	.A(n76));
   NOR4X1M U103 (.Y(N162), 
	.D(n77), 
	.C(n78), 
	.B(n79), 
	.A(n80));
   CLKINVX1M U104 (.Y(o_div_clk), 
	.A(n230));
   OAI211X1M U105 (.Y(next_state[1]), 
	.C0(n124), 
	.B0(n83), 
	.A1(n82), 
	.A0(n81));
   AOI2B1X1M U106 (.Y(n124), 
	.B0(n127), 
	.A1N(n125), 
	.A0(n126));
   AOI21X1M U107 (.Y(n81), 
	.B0(n129), 
	.A1(n128), 
	.A0(n229));
   NAND4X1M U108 (.Y(next_state[0]), 
	.D(n133), 
	.C(n132), 
	.B(n131), 
	.A(n130));
   AOI221XLM U109 (.Y(n133), 
	.C0(n127), 
	.B1(n82), 
	.B0(n134), 
	.A1(n187), 
	.A0(n129));
   OAI2BB1X1M U110 (.Y(n127), 
	.B0(n135), 
	.A1N(N162), 
	.A0N(n134));
   OAI21X1M U111 (.Y(n135), 
	.B0(LTIE_LTIELO_NET), 
	.A1(n136), 
	.A0(n126));
   NOR3X1M U112 (.Y(n129), 
	.C(current_state[0]), 
	.B(current_state[2]), 
	.A(n137));
   NOR4BX1M U113 (.Y(n137), 
	.D(LTIE_LTIELO_NET), 
	.C(HTIE_LTIEHI_NET), 
	.B(LTIE_LTIELO_NET), 
	.AN(n138));
   NOR4X1M U114 (.Y(n138), 
	.D(LTIE_LTIELO_NET), 
	.C(LTIE_LTIELO_NET), 
	.B(LTIE_LTIELO_NET), 
	.A(LTIE_LTIELO_NET));
   NAND2BX1M U115 (.Y(n132), 
	.B(n136), 
	.AN(n139));
   OAI32X1M U116 (.Y(n186), 
	.B1(n141), 
	.B0(n82), 
	.A2(n140), 
	.A1(n187), 
	.A0(n128));
   CLKINVX1M U117 (.Y(n82), 
	.A(LTIE_LTIELO_NET));
   AO22X1M U118 (.Y(n213), 
	.B1(n143), 
	.B0(N28), 
	.A1(Counter_1[3]), 
	.A0(n142));
   AO22X1M U119 (.Y(n214), 
	.B1(n143), 
	.B0(N29), 
	.A1(Counter_1[4]), 
	.A0(n142));
   AO22X1M U120 (.Y(n215), 
	.B1(n143), 
	.B0(N30), 
	.A1(Counter_1[5]), 
	.A0(n142));
   AO22X1M U121 (.Y(n216), 
	.B1(n143), 
	.B0(N31), 
	.A1(Counter_1[6]), 
	.A0(n142));
   AO22X1M U122 (.Y(n217), 
	.B1(n143), 
	.B0(N32), 
	.A1(Counter_1[7]), 
	.A0(n142));
   OAI2BB2X1M U123 (.Y(n218), 
	.B1(n145), 
	.B0(n144), 
	.A1N(n143), 
	.A0N(N33));
   AO22X1M U124 (.Y(n219), 
	.B1(n146), 
	.B0(N36), 
	.A1(n142), 
	.A0(Counter_2[0]));
   AO22X1M U125 (.Y(n220), 
	.B1(n146), 
	.B0(N37), 
	.A1(n142), 
	.A0(Counter_2[1]));
   AO22X1M U126 (.Y(n221), 
	.B1(n146), 
	.B0(N38), 
	.A1(n142), 
	.A0(Counter_2[2]));
   AO22X1M U127 (.Y(n222), 
	.B1(n146), 
	.B0(N39), 
	.A1(n142), 
	.A0(Counter_2[3]));
   AO22X1M U128 (.Y(n223), 
	.B1(n146), 
	.B0(N40), 
	.A1(n142), 
	.A0(Counter_2[4]));
   AO22X1M U129 (.Y(n224), 
	.B1(n146), 
	.B0(N41), 
	.A1(n142), 
	.A0(Counter_2[5]));
   AO22X1M U130 (.Y(n225), 
	.B1(n146), 
	.B0(N42), 
	.A1(n142), 
	.A0(Counter_2[6]));
   AO22X1M U131 (.Y(n226), 
	.B1(n146), 
	.B0(N43), 
	.A1(n142), 
	.A0(Counter_2[7]));
   AO22X1M U132 (.Y(n227), 
	.B1(n146), 
	.B0(N44), 
	.A1(n142), 
	.A0(Counter_2[8]));
   AO22X1M U133 (.Y(n228), 
	.B1(n146), 
	.B0(N45), 
	.A1(n142), 
	.A0(Counter_2[9]));
   OAI2BB2X1M U134 (.Y(n189), 
	.B1(n147), 
	.B0(n144), 
	.A1N(n143), 
	.A0N(N34));
   CLKINVX1M U135 (.Y(n144), 
	.A(n142));
   OAI2BB2X1M U136 (.Y(n190), 
	.B1(n149), 
	.B0(n148), 
	.A1N(n150), 
	.A0N(N56));
   AO2B2X1M U137 (.Y(n191), 
	.B1(n150), 
	.B0(N47), 
	.A1N(n148), 
	.A0(Counter_3[0]));
   AO2B2X1M U138 (.Y(n192), 
	.B1(n150), 
	.B0(N48), 
	.A1N(n2), 
	.A0(Counter_3[1]));
   AO2B2X1M U139 (.Y(n193), 
	.B1(n150), 
	.B0(N49), 
	.A1N(n148), 
	.A0(Counter_3[2]));
   AO2B2X1M U140 (.Y(n194), 
	.B1(n150), 
	.B0(N50), 
	.A1N(n2), 
	.A0(Counter_3[3]));
   AO2B2X1M U141 (.Y(n195), 
	.B1(n150), 
	.B0(N51), 
	.A1N(n148), 
	.A0(Counter_3[4]));
   AO2B2X1M U142 (.Y(n196), 
	.B1(n150), 
	.B0(N52), 
	.A1N(n2), 
	.A0(Counter_3[5]));
   AO2B2X1M U143 (.Y(n197), 
	.B1(n150), 
	.B0(N53), 
	.A1N(n148), 
	.A0(Counter_3[6]));
   AO2B2X1M U144 (.Y(n198), 
	.B1(n150), 
	.B0(N54), 
	.A1N(n2), 
	.A0(Counter_3[7]));
   OAI2BB2X1M U145 (.Y(n199), 
	.B1(n151), 
	.B0(n2), 
	.A1N(n150), 
	.A0N(N55));
   AO2B2X1M U146 (.Y(n200), 
	.B1(n152), 
	.B0(N58), 
	.A1N(n148), 
	.A0(Counter_4[0]));
   AO2B2X1M U147 (.Y(n201), 
	.B1(n152), 
	.B0(N59), 
	.A1N(n2), 
	.A0(Counter_4[1]));
   AO2B2X1M U148 (.Y(n202), 
	.B1(n152), 
	.B0(N60), 
	.A1N(n148), 
	.A0(Counter_4[2]));
   AO2B2X1M U149 (.Y(n203), 
	.B1(n152), 
	.B0(N61), 
	.A1N(n2), 
	.A0(Counter_4[3]));
   AO2B2X1M U150 (.Y(n204), 
	.B1(n152), 
	.B0(N62), 
	.A1N(n148), 
	.A0(Counter_4[4]));
   AO2B2X1M U151 (.Y(n205), 
	.B1(n152), 
	.B0(N63), 
	.A1N(n2), 
	.A0(Counter_4[5]));
   AO2B2X1M U152 (.Y(n206), 
	.B1(n152), 
	.B0(N64), 
	.A1N(n148), 
	.A0(Counter_4[6]));
   AO2B2X1M U153 (.Y(n207), 
	.B1(n152), 
	.B0(N65), 
	.A1N(n2), 
	.A0(Counter_4[7]));
   OAI2BB2X1M U154 (.Y(n208), 
	.B1(n153), 
	.B0(n148), 
	.A1N(n152), 
	.A0N(N66));
   OAI2BB2X1M U155 (.Y(n209), 
	.B1(n154), 
	.B0(n2), 
	.A1N(n152), 
	.A0N(N67));
   NAND2BX1M U156 (.Y(n141), 
	.B(n134), 
	.AN(N162));
   NOR3X1M U157 (.Y(n134), 
	.C(n188), 
	.B(current_state[1]), 
	.A(current_state[0]));
   AO22X1M U158 (.Y(n210), 
	.B1(n143), 
	.B0(N25), 
	.A1(Counter_1[0]), 
	.A0(n142));
   AO22X1M U159 (.Y(n211), 
	.B1(n143), 
	.B0(N26), 
	.A1(Counter_1[1]), 
	.A0(n142));
   AO22X1M U160 (.Y(n212), 
	.B1(n143), 
	.B0(N27), 
	.A1(Counter_1[2]), 
	.A0(n142));
   NAND3X1M U161 (.Y(n130), 
	.C(n229), 
	.B(current_state[1]), 
	.A(n128));
   CLKINVX1M U162 (.Y(n229), 
	.A(n140));
   NAND4X1M U163 (.Y(n128), 
	.D(n158), 
	.C(n157), 
	.B(n156), 
	.A(n155));
   NOR4X1M U164 (.Y(n158), 
	.D(n161), 
	.C(Counter_1[7]), 
	.B(n160), 
	.A(n159));
   CLKXOR2X2M U165 (.Y(n161), 
	.B(Counter_1[0]), 
	.A(even_ratio[0]));
   CLKXOR2X2M U166 (.Y(n160), 
	.B(Counter_1[5]), 
	.A(even_ratio[5]));
   NAND3X1M U167 (.Y(n159), 
	.C(n145), 
	.B(n162), 
	.A(n147));
   CLKINVX1M U168 (.Y(n145), 
	.A(Counter_1[8]));
   CLKINVX1M U169 (.Y(n147), 
	.A(Counter_1[9]));
   NOR3X1M U170 (.Y(n157), 
	.C(n165), 
	.B(n164), 
	.A(n163));
   CLKXOR2X2M U171 (.Y(n165), 
	.B(Counter_1[1]), 
	.A(even_ratio[1]));
   CLKXOR2X2M U172 (.Y(n164), 
	.B(Counter_1[3]), 
	.A(even_ratio[3]));
   CLKXOR2X2M U173 (.Y(n163), 
	.B(Counter_1[2]), 
	.A(even_ratio[2]));
   XNOR2X1M U174 (.Y(n156), 
	.B(even_ratio[4]), 
	.A(Counter_1[4]));
   XNOR2X1M U175 (.Y(n155), 
	.B(even_ratio[6]), 
	.A(Counter_1[6]));
   CLKNAND2X2M U176 (.Y(n131), 
	.B(n125), 
	.A(n126));
   NAND4X1M U177 (.Y(n125), 
	.D(n169), 
	.C(n168), 
	.B(n167), 
	.A(n166));
   NOR4X1M U178 (.Y(n169), 
	.D(n172), 
	.C(Counter_3[7]), 
	.B(n171), 
	.A(n170));
   CLKXOR2X2M U179 (.Y(n172), 
	.B(Counter_3[0]), 
	.A(even_ratio[0]));
   CLKXOR2X2M U180 (.Y(n171), 
	.B(Counter_3[5]), 
	.A(even_ratio[5]));
   NAND3X1M U181 (.Y(n170), 
	.C(n151), 
	.B(n162), 
	.A(n149));
   CLKINVX1M U182 (.Y(n151), 
	.A(Counter_3[8]));
   CLKINVX1M U183 (.Y(n149), 
	.A(Counter_3[9]));
   NOR3X1M U184 (.Y(n168), 
	.C(n175), 
	.B(n174), 
	.A(n173));
   CLKXOR2X2M U185 (.Y(n175), 
	.B(Counter_3[1]), 
	.A(even_ratio[1]));
   CLKXOR2X2M U186 (.Y(n174), 
	.B(Counter_3[3]), 
	.A(even_ratio[3]));
   CLKXOR2X2M U187 (.Y(n173), 
	.B(Counter_3[2]), 
	.A(even_ratio[2]));
   XNOR2X1M U188 (.Y(n167), 
	.B(even_ratio[4]), 
	.A(Counter_3[4]));
   XNOR2X1M U189 (.Y(n166), 
	.B(even_ratio[6]), 
	.A(Counter_3[6]));
   NOR2X1M U190 (.Y(n126), 
	.B(current_state[1]), 
	.A(n140));
   CLKNAND2X2M U191 (.Y(n140), 
	.B(n188), 
	.A(current_state[0]));
   CLKINVX1M U192 (.Y(n188), 
	.A(current_state[2]));
   CLKNAND2X2M U193 (.Y(n83), 
	.B(n139), 
	.A(n136));
   NAND4X1M U194 (.Y(n139), 
	.D(n179), 
	.C(n178), 
	.B(n177), 
	.A(n176));
   NOR4X1M U195 (.Y(n179), 
	.D(n182), 
	.C(Counter_4[7]), 
	.B(n181), 
	.A(n180));
   CLKXOR2X2M U196 (.Y(n182), 
	.B(Counter_4[0]), 
	.A(even_ratio[0]));
   CLKXOR2X2M U197 (.Y(n181), 
	.B(Counter_4[5]), 
	.A(even_ratio[5]));
   NAND3X1M U198 (.Y(n180), 
	.C(n153), 
	.B(n162), 
	.A(n154));
   CLKINVX1M U199 (.Y(n153), 
	.A(Counter_4[8]));
   CLKINVX1M U200 (.Y(n162), 
	.A(even_ratio_31));
   CLKINVX1M U201 (.Y(n154), 
	.A(Counter_4[9]));
   NOR3X1M U202 (.Y(n178), 
	.C(n185), 
	.B(n184), 
	.A(n183));
   CLKXOR2X2M U203 (.Y(n185), 
	.B(Counter_4[1]), 
	.A(even_ratio[1]));
   CLKXOR2X2M U204 (.Y(n184), 
	.B(Counter_4[3]), 
	.A(even_ratio[3]));
   CLKXOR2X2M U205 (.Y(n183), 
	.B(Counter_4[2]), 
	.A(even_ratio[2]));
   XNOR2X1M U206 (.Y(n177), 
	.B(even_ratio[4]), 
	.A(Counter_4[4]));
   XNOR2X1M U207 (.Y(n176), 
	.B(even_ratio[6]), 
	.A(Counter_4[6]));
   NOR3X1M U208 (.Y(n136), 
	.C(n187), 
	.B(current_state[2]), 
	.A(current_state[0]));
   CLKINVX1M U209 (.Y(n187), 
	.A(current_state[1]));
   ClkDiv___1_DW01_inc_0 add_72 (.A({ Counter_4[9],
		Counter_4[8],
		Counter_4[7],
		Counter_4[6],
		Counter_4[5],
		Counter_4[4],
		Counter_4[3],
		Counter_4[2],
		Counter_4[1],
		Counter_4[0] }), 
	.SUM({ N67,
		N66,
		N65,
		N64,
		N63,
		N62,
		N61,
		N60,
		N59,
		N58 }));
   ClkDiv___1_DW01_inc_1 add_67 (.A({ Counter_3[9],
		Counter_3[8],
		Counter_3[7],
		Counter_3[6],
		Counter_3[5],
		Counter_3[4],
		Counter_3[3],
		Counter_3[2],
		Counter_3[1],
		Counter_3[0] }), 
	.SUM({ N56,
		N55,
		N54,
		N53,
		N52,
		N51,
		N50,
		N49,
		N48,
		N47 }));
   ClkDiv___1_DW01_inc_2 add_62 (.A({ Counter_2[9],
		Counter_2[8],
		Counter_2[7],
		Counter_2[6],
		Counter_2[5],
		Counter_2[4],
		Counter_2[3],
		Counter_2[2],
		Counter_2[1],
		Counter_2[0] }), 
	.SUM({ N45,
		N44,
		N43,
		N42,
		N41,
		N40,
		N39,
		N38,
		N37,
		N36 }));
   ClkDiv___1_DW01_inc_3 add_57 (.A({ Counter_1[9],
		Counter_1[8],
		Counter_1[7],
		Counter_1[6],
		Counter_1[5],
		Counter_1[4],
		Counter_1[3],
		Counter_1[2],
		Counter_1[1],
		Counter_1[0] }), 
	.SUM({ N34,
		N33,
		N32,
		N31,
		N30,
		N29,
		N28,
		N27,
		N26,
		N25 }));
   NAND3BX2M U3 (.Y(n79), 
	.C(n68), 
	.B(n67), 
	.AN(n80));
endmodule

module Rst_Sync_NUM_STAGES2_ACTIVE_TYPLOW_test_0 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_so, 
	test_se);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   output test_so;
   input test_se;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [1:0] FF_Stage;

   assign test_so = FF_Stage[1] ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRQX2M \FF_Stage_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(RST), 
	.Q(FF_Stage[0]), 
	.D(HTIE_LTIEHI_NET), 
	.CK(CLK));
   SDFFRQX1M \FF_Stage_reg[1]  (.SI(FF_Stage[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(FF_Stage[1]), 
	.D(FF_Stage[0]), 
	.CK(CLK));
   AND2X2M U6 (.Y(SYNC_RST), 
	.B(RST), 
	.A(FF_Stage[1]));
endmodule

module Rst_Sync_NUM_STAGES2_ACTIVE_TYPLOW_test_1 (
	RST, 
	CLK, 
	SYNC_RST, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN22_SE);
   input RST;
   input CLK;
   output SYNC_RST;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN22_SE;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [1:0] FF_Stage;

   assign test_so = FF_Stage[1] ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRQX2M \FF_Stage_reg[0]  (.SI(test_si), 
	.SE(FE_OFN22_SE), 
	.RN(RST), 
	.Q(FF_Stage[0]), 
	.D(HTIE_LTIEHI_NET), 
	.CK(CLK));
   SDFFRQX1M \FF_Stage_reg[1]  (.SI(FF_Stage[0]), 
	.SE(test_se), 
	.RN(RST), 
	.Q(FF_Stage[1]), 
	.D(FF_Stage[0]), 
	.CK(CLK));
   AND2X2M U6 (.Y(SYNC_RST), 
	.B(RST), 
	.A(FF_Stage[1]));
endmodule

module Data_Sync_NUM_STAGES2_BUS_WIDTH8_test_1 (
	CLK, 
	RST_n, 
	bus_enable, 
	UNSYNC_bus, 
	enable_pulse, 
	SYNC_bus, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN8_RST_D1_M, 
	FE_OFN18_SE, 
	REF_CLK_M__L5_N1);
   input CLK;
   input RST_n;
   input bus_enable;
   input [7:0] UNSYNC_bus;
   output enable_pulse;
   output [7:0] SYNC_bus;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN8_RST_D1_M;
   input FE_OFN18_SE;
   input REF_CLK_M__L5_N1;

   // Internal wires
   wire pulse_gen;
   wire Q_in;
   wire N3;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n19;
   wire n1;
   wire n2;
   wire [1:0] FF_Stage;

   assign test_so2 = pulse_gen ;
   assign test_so1 = Q_in ;

   SDFFRQX2M \FF_Stage_reg[1]  (.SI(FF_Stage[0]), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(FF_Stage[1]), 
	.D(FF_Stage[0]), 
	.CK(CLK));
   SDFFRQX2M Q_in_reg (.SI(FF_Stage[1]), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(Q_in), 
	.D(FF_Stage[1]), 
	.CK(CLK));
   SDFFRQX2M \SYNC_bus_reg[7]  (.SI(SYNC_bus[6]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[7]), 
	.D(n19), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \SYNC_bus_reg[4]  (.SI(SYNC_bus[3]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[4]), 
	.D(n13), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \SYNC_bus_reg[6]  (.SI(SYNC_bus[5]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[6]), 
	.D(n17), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \SYNC_bus_reg[5]  (.SI(SYNC_bus[4]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[5]), 
	.D(n15), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M pulse_gen_reg (.SI(enable_pulse), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(pulse_gen), 
	.D(N3), 
	.CK(CLK));
   SDFFRQX2M \SYNC_bus_reg[3]  (.SI(SYNC_bus[2]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[3]), 
	.D(n11), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \SYNC_bus_reg[0]  (.SI(test_si2), 
	.SE(test_se), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[0]), 
	.D(n5), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \SYNC_bus_reg[2]  (.SI(SYNC_bus[1]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[2]), 
	.D(n9), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \SYNC_bus_reg[1]  (.SI(SYNC_bus[0]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(SYNC_bus[1]), 
	.D(n7), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M enable_pulse_reg (.SI(SYNC_bus[7]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(enable_pulse), 
	.D(pulse_gen), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0]  (.SI(test_si1), 
	.SE(test_se), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(FF_Stage[0]), 
	.D(bus_enable), 
	.CK(CLK));
   AO22X1M U3 (.Y(n5), 
	.B1(n2), 
	.B0(SYNC_bus[0]), 
	.A1(UNSYNC_bus[0]), 
	.A0(pulse_gen));
   AO22X1M U4 (.Y(n7), 
	.B1(n2), 
	.B0(SYNC_bus[1]), 
	.A1(pulse_gen), 
	.A0(UNSYNC_bus[1]));
   AO22X1M U5 (.Y(n9), 
	.B1(n2), 
	.B0(SYNC_bus[2]), 
	.A1(pulse_gen), 
	.A0(UNSYNC_bus[2]));
   AO22X1M U6 (.Y(n11), 
	.B1(n2), 
	.B0(SYNC_bus[3]), 
	.A1(pulse_gen), 
	.A0(UNSYNC_bus[3]));
   AO22X1M U7 (.Y(n13), 
	.B1(n2), 
	.B0(SYNC_bus[4]), 
	.A1(pulse_gen), 
	.A0(UNSYNC_bus[4]));
   AO22X1M U8 (.Y(n15), 
	.B1(n2), 
	.B0(SYNC_bus[5]), 
	.A1(pulse_gen), 
	.A0(UNSYNC_bus[5]));
   AO22X1M U9 (.Y(n17), 
	.B1(n2), 
	.B0(SYNC_bus[6]), 
	.A1(pulse_gen), 
	.A0(UNSYNC_bus[6]));
   AO22X1M U10 (.Y(n19), 
	.B1(n2), 
	.B0(SYNC_bus[7]), 
	.A1(pulse_gen), 
	.A0(UNSYNC_bus[7]));
   INVX2M U11 (.Y(n2), 
	.A(pulse_gen));
   AND3X2M U12 (.Y(N3), 
	.C(FE_OFN8_RST_D1_M), 
	.B(FF_Stage[1]), 
	.A(n1));
   INVX2M U13 (.Y(n1), 
	.A(Q_in));
endmodule

module SYS_CTRL_test_1 (
	CLK, 
	RST, 
	Data_sync, 
	enable_pulse, 
	FIFO_FULL, 
	Rd_DATA, 
	Rd_Valid, 
	ALU_OUT, 
	OUT_VALID, 
	WR_DATA, 
	WR_INC, 
	FUN, 
	EN, 
	Gate_En, 
	Wr_D, 
	Addr, 
	RdEn, 
	WrEn, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN11_RST_D1_M, 
	FE_OFN12_RST_D1_M, 
	FE_OFN8_RST_D1_M, 
	FE_OFN18_SE, 
	FE_OFN19_SE, 
	REF_CLK_M__L5_N1, 
	REF_CLK_M__L5_N2);
   input CLK;
   input RST;
   input [7:0] Data_sync;
   input enable_pulse;
   input FIFO_FULL;
   input [7:0] Rd_DATA;
   input Rd_Valid;
   input [15:0] ALU_OUT;
   input OUT_VALID;
   output [7:0] WR_DATA;
   output WR_INC;
   output [3:0] FUN;
   output EN;
   output Gate_En;
   output [7:0] Wr_D;
   output [7:0] Addr;
   output RdEn;
   output WrEn;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN11_RST_D1_M;
   input FE_OFN12_RST_D1_M;
   input FE_OFN8_RST_D1_M;
   input FE_OFN18_SE;
   input FE_OFN19_SE;
   input REF_CLK_M__L5_N1;
   input REF_CLK_M__L5_N2;

   // Internal wires
   wire FE_OFN16_Addr_2_;
   wire flag_1;
   wire N225;
   wire N226;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n92;
   wire [3:0] current_state;
   wire [3:0] next_state;
   wire [1:0] Counter;
   wire [7:0] Addr_next;

   assign test_so = flag_1 ;

   BUFX2M FE_OFC16_Addr_2_ (.Y(Addr[2]), 
	.A(FE_OFN16_Addr_2_));
   SDFFRQX2M \Addr_next_reg[7]  (.SI(Addr_next[6]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[7]), 
	.D(Addr[7]), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \Addr_next_reg[6]  (.SI(Addr_next[5]), 
	.SE(test_se), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[6]), 
	.D(Addr[6]), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \Addr_next_reg[5]  (.SI(Addr_next[4]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[5]), 
	.D(Addr[5]), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \Addr_next_reg[4]  (.SI(Addr_next[3]), 
	.SE(test_se), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[4]), 
	.D(Addr[4]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Addr_next_reg[3]  (.SI(Addr_next[2]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[3]), 
	.D(Addr[3]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Addr_next_reg[2]  (.SI(Addr_next[1]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[2]), 
	.D(Addr[2]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Addr_next_reg[1]  (.SI(Addr_next[0]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[1]), 
	.D(Addr[1]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Addr_next_reg[0]  (.SI(test_si), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Addr_next[0]), 
	.D(Addr[0]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M flag_1_reg (.SI(current_state[3]), 
	.SE(test_se), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(flag_1), 
	.D(n19), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Counter_reg[1]  (.SI(Counter[0]), 
	.SE(FE_OFN18_SE), 
	.RN(RST), 
	.Q(Counter[1]), 
	.D(N226), 
	.CK(CLK));
   SDFFRQX2M \Counter_reg[0]  (.SI(Addr_next[7]), 
	.SE(test_se), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(Counter[0]), 
	.D(N225), 
	.CK(REF_CLK_M__L5_N1));
   SDFFRQX2M \current_state_reg[2]  (.SI(current_state[1]), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(current_state[2]), 
	.D(next_state[2]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \current_state_reg[3]  (.SI(current_state[2]), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(current_state[3]), 
	.D(next_state[3]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \current_state_reg[0]  (.SI(Counter[1]), 
	.SE(test_se), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \current_state_reg[1]  (.SI(n28), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(current_state[1]), 
	.D(next_state[1]), 
	.CK(REF_CLK_M__L5_N2));
   NOR2X2M U18 (.Y(FUN[3]), 
	.B(n33), 
	.A(n17));
   NOR2X2M U19 (.Y(FUN[1]), 
	.B(n35), 
	.A(n17));
   INVX2M U21 (.Y(n92), 
	.A(enable_pulse));
   OAI21X2M U22 (.Y(FE_OFN16_Addr_2_), 
	.B0(n88), 
	.A1(n34), 
	.A0(n80));
   OAI21X2M U23 (.Y(EN), 
	.B0(n38), 
	.A1(n37), 
	.A0(OUT_VALID));
   INVX2M U24 (.Y(n23), 
	.A(n57));
   NAND2X2M U25 (.Y(n83), 
	.B(n52), 
	.A(n61));
   INVX2M U26 (.Y(n21), 
	.A(n91));
   INVX2M U27 (.Y(n22), 
	.A(n43));
   NOR2BX2M U28 (.Y(Wr_D[0]), 
	.B(n65), 
	.AN(n72));
   NOR2BX2M U29 (.Y(Wr_D[1]), 
	.B(n65), 
	.AN(n71));
   NOR2BX2M U30 (.Y(Wr_D[2]), 
	.B(n65), 
	.AN(n70));
   NOR2BX2M U31 (.Y(Wr_D[3]), 
	.B(n65), 
	.AN(n69));
   NOR2BX2M U32 (.Y(Wr_D[4]), 
	.B(n65), 
	.AN(n68));
   NOR2BX2M U33 (.Y(Wr_D[5]), 
	.B(n65), 
	.AN(n67));
   NOR2BX2M U34 (.Y(Wr_D[6]), 
	.B(n65), 
	.AN(n66));
   NOR2X2M U35 (.Y(n57), 
	.B(n75), 
	.A(n74));
   NAND2X2M U36 (.Y(n55), 
	.B(n46), 
	.A(n61));
   AOI21X2M U37 (.Y(n80), 
	.B0(n47), 
	.A1(n21), 
	.A0(n92));
   NOR2X2M U38 (.Y(n82), 
	.B(n92), 
	.A(n91));
   NOR2X2M U39 (.Y(FUN[2]), 
	.B(n34), 
	.A(n17));
   NAND2X2M U40 (.Y(n52), 
	.B(n27), 
	.A(n62));
   NAND3X2M U41 (.Y(n37), 
	.C(n40), 
	.B(n24), 
	.A(n28));
   NAND2X2M U42 (.Y(n42), 
	.B(n73), 
	.A(n27));
   NAND2X2M U43 (.Y(n61), 
	.B(n76), 
	.A(n62));
   NOR2X3M U44 (.Y(FUN[0]), 
	.B(n36), 
	.A(n17));
   NAND2X2M U45 (.Y(n91), 
	.B(n77), 
	.A(n62));
   INVX2M U46 (.Y(n17), 
	.A(Gate_En));
   NAND2X2M U47 (.Y(n46), 
	.B(n73), 
	.A(n76));
   NOR2X2M U48 (.Y(n72), 
	.B(n92), 
	.A(n36));
   NAND2X2M U49 (.Y(n43), 
	.B(n77), 
	.A(n73));
   NOR2X2M U50 (.Y(WR_INC), 
	.B(n57), 
	.A(FIFO_FULL));
   INVX2M U51 (.Y(n19), 
	.A(n79));
   INVX2M U52 (.Y(n27), 
	.A(n41));
   NOR2X2M U53 (.Y(Wr_D[7]), 
	.B(n64), 
	.A(n65));
   OAI21X2M U54 (.Y(RdEn), 
	.B0(n18), 
	.A1(n52), 
	.A0(n92));
   NOR3BX4M U55 (.Y(n65), 
	.C(n21), 
	.B(n48), 
	.AN(n46));
   AND2X2M U56 (.Y(n74), 
	.B(n77), 
	.A(n40));
   AND2X2M U57 (.Y(n75), 
	.B(n40), 
	.A(n76));
   NOR2X2M U58 (.Y(n71), 
	.B(n92), 
	.A(n35));
   NOR2X2M U59 (.Y(n70), 
	.B(n92), 
	.A(n34));
   NOR2X2M U60 (.Y(n69), 
	.B(n92), 
	.A(n33));
   INVX2M U61 (.Y(n18), 
	.A(n47));
   NOR2X2M U62 (.Y(WrEn), 
	.B(n92), 
	.A(n65));
   AND4X2M U63 (.Y(n51), 
	.D(n63), 
	.C(n62), 
	.B(n24), 
	.A(n28));
   NOR2X2M U64 (.Y(n63), 
	.B(n33), 
	.A(n64));
   NOR2X2M U65 (.Y(n68), 
	.B(n92), 
	.A(n32));
   NOR2X2M U66 (.Y(n67), 
	.B(n92), 
	.A(n31));
   NOR2X2M U67 (.Y(n66), 
	.B(n92), 
	.A(n30));
   OAI21X4M U68 (.Y(Addr[3]), 
	.B0(n87), 
	.A1(n33), 
	.A0(n80));
   AOI22X1M U69 (.Y(n87), 
	.B1(n83), 
	.B0(n69), 
	.A1(n82), 
	.A0(Addr_next[3]));
   AOI22X1M U70 (.Y(n88), 
	.B1(n83), 
	.B0(n70), 
	.A1(n82), 
	.A0(Addr_next[2]));
   OAI221X1M U71 (.Y(Addr[0]), 
	.C0(n90), 
	.B1(n46), 
	.B0(n92), 
	.A1(n36), 
	.A0(n80));
   AOI22X1M U72 (.Y(n90), 
	.B1(n83), 
	.B0(n72), 
	.A1(n82), 
	.A0(Addr_next[0]));
   NOR2X2M U73 (.Y(n62), 
	.B(current_state[2]), 
	.A(current_state[3]));
   NOR2BX2M U74 (.Y(n73), 
	.B(current_state[3]), 
	.AN(current_state[2]));
   OAI21X2M U75 (.Y(n79), 
	.B0(n22), 
	.A1(flag_1), 
	.A0(enable_pulse));
   OAI21X2M U76 (.Y(Gate_En), 
	.B0(n79), 
	.A1(n37), 
	.A0(OUT_VALID));
   NOR2X2M U77 (.Y(n77), 
	.B(current_state[0]), 
	.A(n24));
   NOR2X2M U78 (.Y(n76), 
	.B(current_state[1]), 
	.A(n28));
   NOR2BX2M U79 (.Y(n40), 
	.B(current_state[2]), 
	.AN(current_state[3]));
   OAI21X2M U80 (.Y(Addr[1]), 
	.B0(n89), 
	.A1(n35), 
	.A0(n80));
   AOI22X1M U81 (.Y(n89), 
	.B1(n83), 
	.B0(n71), 
	.A1(n82), 
	.A0(Addr_next[1]));
   NOR2X2M U82 (.Y(n47), 
	.B(Rd_Valid), 
	.A(n42));
   AO22X1M U83 (.Y(WR_DATA[0]), 
	.B1(n75), 
	.B0(ALU_OUT[0]), 
	.A1(n74), 
	.A0(Rd_DATA[0]));
   AO22X1M U84 (.Y(WR_DATA[1]), 
	.B1(n75), 
	.B0(ALU_OUT[1]), 
	.A1(n74), 
	.A0(Rd_DATA[1]));
   AO22X1M U85 (.Y(WR_DATA[2]), 
	.B1(n75), 
	.B0(ALU_OUT[2]), 
	.A1(n74), 
	.A0(Rd_DATA[2]));
   AO22X1M U86 (.Y(WR_DATA[3]), 
	.B1(n75), 
	.B0(ALU_OUT[3]), 
	.A1(n74), 
	.A0(Rd_DATA[3]));
   AO22X1M U87 (.Y(WR_DATA[4]), 
	.B1(n75), 
	.B0(ALU_OUT[4]), 
	.A1(n74), 
	.A0(Rd_DATA[4]));
   AO22X1M U88 (.Y(WR_DATA[5]), 
	.B1(n75), 
	.B0(ALU_OUT[5]), 
	.A1(n74), 
	.A0(Rd_DATA[5]));
   AO22X1M U89 (.Y(WR_DATA[6]), 
	.B1(n75), 
	.B0(ALU_OUT[6]), 
	.A1(n74), 
	.A0(Rd_DATA[6]));
   AO22X1M U90 (.Y(WR_DATA[7]), 
	.B1(n75), 
	.B0(ALU_OUT[7]), 
	.A1(n74), 
	.A0(Rd_DATA[7]));
   NAND3X2M U91 (.Y(n38), 
	.C(Counter[1]), 
	.B(n19), 
	.A(Counter[0]));
   NAND2X2M U92 (.Y(n41), 
	.B(current_state[1]), 
	.A(current_state[0]));
   INVX2M U93 (.Y(n28), 
	.A(current_state[0]));
   INVX2M U94 (.Y(n24), 
	.A(current_state[1]));
   NOR3BX2M U95 (.Y(n48), 
	.C(current_state[1]), 
	.B(current_state[0]), 
	.AN(n73));
   NAND3X2M U96 (.Y(next_state[3]), 
	.C(n39), 
	.B(n38), 
	.A(n37));
   AOI32X1M U97 (.Y(n39), 
	.B1(n26), 
	.B0(Rd_Valid), 
	.A2(FIFO_FULL), 
	.A1(n41), 
	.A0(n40));
   INVX2M U98 (.Y(n26), 
	.A(n42));
   INVX2M U99 (.Y(n35), 
	.A(Data_sync[1]));
   INVX2M U100 (.Y(n34), 
	.A(Data_sync[2]));
   NAND4X2M U101 (.Y(next_state[1]), 
	.D(n54), 
	.C(n53), 
	.B(n42), 
	.A(n52));
   AOI222X1M U102 (.Y(n54), 
	.C1(n38), 
	.C0(n22), 
	.B1(n55), 
	.B0(enable_pulse), 
	.A1(n92), 
	.A0(n21));
   AOI32X1M U103 (.Y(n53), 
	.B1(n23), 
	.B0(FIFO_FULL), 
	.A2(n56), 
	.A1(Data_sync[0]), 
	.A0(n51));
   AOI2BB1X2M U104 (.Y(n56), 
	.B0(n32), 
	.A1N(n58), 
	.A0N(n50));
   INVX2M U105 (.Y(n33), 
	.A(Data_sync[3]));
   INVX2M U106 (.Y(n36), 
	.A(Data_sync[0]));
   NOR4X1M U107 (.Y(n58), 
	.D(Data_sync[6]), 
	.C(Data_sync[2]), 
	.B(n35), 
	.A(n31));
   NOR4X1M U108 (.Y(n50), 
	.D(Data_sync[5]), 
	.C(Data_sync[1]), 
	.B(n34), 
	.A(n30));
   OAI2B11X2M U109 (.Y(next_state[2]), 
	.C0(n45), 
	.B0(n44), 
	.A1N(n38), 
	.A0(n43));
   AOI32X1M U110 (.Y(n44), 
	.B1(Rd_Valid), 
	.B0(n25), 
	.A2(n51), 
	.A1(n50), 
	.A0(n49));
   NOR3BX2M U111 (.Y(n45), 
	.C(n48), 
	.B(n47), 
	.AN(n46));
   INVX2M U112 (.Y(n25), 
	.A(n52));
   NAND2X2M U113 (.Y(n64), 
	.B(Data_sync[7]), 
	.A(enable_pulse));
   OAI2B1X2M U114 (.Y(Addr[7]), 
	.B0(n81), 
	.A1N(Data_sync[7]), 
	.A0(n80));
   AOI22X1M U115 (.Y(n81), 
	.B1(n83), 
	.B0(n29), 
	.A1(n82), 
	.A0(Addr_next[7]));
   INVX2M U116 (.Y(n29), 
	.A(n64));
   OAI21X2M U117 (.Y(Addr[4]), 
	.B0(n86), 
	.A1(n32), 
	.A0(n80));
   AOI22X1M U118 (.Y(n86), 
	.B1(n83), 
	.B0(n68), 
	.A1(n82), 
	.A0(Addr_next[4]));
   OAI21X2M U119 (.Y(Addr[5]), 
	.B0(n85), 
	.A1(n31), 
	.A0(n80));
   AOI22X1M U120 (.Y(n85), 
	.B1(n83), 
	.B0(n67), 
	.A1(n82), 
	.A0(Addr_next[5]));
   OAI21X2M U121 (.Y(Addr[6]), 
	.B0(n84), 
	.A1(n30), 
	.A0(n80));
   AOI22X1M U122 (.Y(n84), 
	.B1(n83), 
	.B0(n66), 
	.A1(n82), 
	.A0(Addr_next[6]));
   NOR2X2M U123 (.Y(N225), 
	.B(enable_pulse), 
	.A(Counter[0]));
   NAND4X2M U124 (.Y(next_state[0]), 
	.D(n60), 
	.C(n59), 
	.B(n18), 
	.A(n52));
   NAND3X2M U125 (.Y(n59), 
	.C(n58), 
	.B(n51), 
	.A(n49));
   AOI222X1M U126 (.Y(n60), 
	.C1(n20), 
	.C0(OUT_VALID), 
	.B1(n92), 
	.B0(n55), 
	.A1(enable_pulse), 
	.A0(n48));
   INVX2M U127 (.Y(n20), 
	.A(n37));
   INVX2M U128 (.Y(n31), 
	.A(Data_sync[5]));
   INVX2M U129 (.Y(n30), 
	.A(Data_sync[6]));
   AOI2BB1X2M U130 (.Y(N226), 
	.B0(n78), 
	.A1N(Counter[1]), 
	.A0N(Counter[0]));
   AOI2B1X1M U131 (.Y(n78), 
	.B0(N225), 
	.A1N(Counter[1]), 
	.A0(n92));
   INVX2M U132 (.Y(n32), 
	.A(Data_sync[4]));
   CLKXOR2X2M U133 (.Y(n49), 
	.B(Data_sync[4]), 
	.A(n36));
endmodule

module Register_File_10_0_1_test_1 (
	CLK, 
	RST_n, 
	RdEn, 
	WrEn, 
	Address, 
	WrData, 
	RdData, 
	RdData_Valid, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN10_RST_D1_M, 
	FE_OFN11_RST_D1_M, 
	FE_OFN8_RST_D1_M, 
	FE_OFN18_SE, 
	FE_OFN19_SE, 
	FE_OFN22_SE, 
	REF_CLK_M__L5_N2, 
	REF_CLK_M__L5_N5, 
	REF_CLK_M__L5_N6);
   input CLK;
   input RST_n;
   input RdEn;
   input WrEn;
   input [3:0] Address;
   input [7:0] WrData;
   output [7:0] RdData;
   output RdData_Valid;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN10_RST_D1_M;
   input FE_OFN11_RST_D1_M;
   input FE_OFN8_RST_D1_M;
   input FE_OFN18_SE;
   input FE_OFN19_SE;
   input FE_OFN22_SE;
   input REF_CLK_M__L5_N2;
   input REF_CLK_M__L5_N5;
   input REF_CLK_M__L5_N6;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire FE_OFN33_REG0_2_;
   wire FE_OFN32_REG0_3_;
   wire FE_OFN31_REG0_4_;
   wire FE_OFN30_REG0_5_;
   wire FE_OFN29_REG0_6_;
   wire FE_OFN28_REG0_7_;
   wire FE_OFN27_REG1_7_;
   wire FE_OFN26_REG1_6_;
   wire FE_OFN25_SE;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire \reg_file[4][7] ;
   wire \reg_file[4][6] ;
   wire \reg_file[4][5] ;
   wire \reg_file[4][4] ;
   wire \reg_file[4][3] ;
   wire \reg_file[4][2] ;
   wire \reg_file[4][1] ;
   wire \reg_file[4][0] ;
   wire \reg_file[5][7] ;
   wire \reg_file[5][6] ;
   wire \reg_file[5][5] ;
   wire \reg_file[5][4] ;
   wire \reg_file[5][3] ;
   wire \reg_file[5][2] ;
   wire \reg_file[5][1] ;
   wire \reg_file[5][0] ;
   wire \reg_file[6][7] ;
   wire \reg_file[6][6] ;
   wire \reg_file[6][5] ;
   wire \reg_file[6][4] ;
   wire \reg_file[6][3] ;
   wire \reg_file[6][2] ;
   wire \reg_file[6][1] ;
   wire \reg_file[6][0] ;
   wire \reg_file[7][7] ;
   wire \reg_file[7][6] ;
   wire \reg_file[7][5] ;
   wire \reg_file[7][4] ;
   wire \reg_file[7][3] ;
   wire \reg_file[7][2] ;
   wire \reg_file[7][1] ;
   wire \reg_file[7][0] ;
   wire \reg_file[8][7] ;
   wire \reg_file[8][6] ;
   wire \reg_file[8][5] ;
   wire \reg_file[8][4] ;
   wire \reg_file[8][3] ;
   wire \reg_file[8][2] ;
   wire \reg_file[8][1] ;
   wire \reg_file[8][0] ;
   wire \reg_file[9][7] ;
   wire \reg_file[9][6] ;
   wire \reg_file[9][5] ;
   wire \reg_file[9][4] ;
   wire \reg_file[9][3] ;
   wire \reg_file[9][2] ;
   wire \reg_file[9][1] ;
   wire \reg_file[9][0] ;
   wire \reg_file[10][7] ;
   wire \reg_file[10][6] ;
   wire \reg_file[10][5] ;
   wire \reg_file[10][4] ;
   wire \reg_file[10][3] ;
   wire \reg_file[10][2] ;
   wire \reg_file[10][1] ;
   wire \reg_file[10][0] ;
   wire \reg_file[11][7] ;
   wire \reg_file[11][6] ;
   wire \reg_file[11][5] ;
   wire \reg_file[11][4] ;
   wire \reg_file[11][3] ;
   wire \reg_file[11][2] ;
   wire \reg_file[11][1] ;
   wire \reg_file[11][0] ;
   wire \reg_file[12][7] ;
   wire \reg_file[12][6] ;
   wire \reg_file[12][5] ;
   wire \reg_file[12][4] ;
   wire \reg_file[12][3] ;
   wire \reg_file[12][2] ;
   wire \reg_file[12][1] ;
   wire \reg_file[12][0] ;
   wire \reg_file[13][7] ;
   wire \reg_file[13][6] ;
   wire \reg_file[13][5] ;
   wire \reg_file[13][4] ;
   wire \reg_file[13][3] ;
   wire \reg_file[13][2] ;
   wire \reg_file[13][1] ;
   wire \reg_file[13][0] ;
   wire \reg_file[14][7] ;
   wire \reg_file[14][6] ;
   wire \reg_file[14][5] ;
   wire \reg_file[14][4] ;
   wire \reg_file[14][3] ;
   wire \reg_file[14][2] ;
   wire \reg_file[14][1] ;
   wire \reg_file[14][0] ;
   wire \reg_file[15][7] ;
   wire \reg_file[15][6] ;
   wire \reg_file[15][5] ;
   wire \reg_file[15][4] ;
   wire \reg_file[15][3] ;
   wire \reg_file[15][2] ;
   wire \reg_file[15][1] ;
   wire \reg_file[15][0] ;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n357;
   wire n358;
   wire n359;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;

   assign N10 = Address[0] ;
   assign N11 = Address[1] ;
   assign N12 = Address[2] ;
   assign N13 = Address[3] ;
   assign test_so1 = \reg_file[11][4]  ;
   assign test_so2 = \reg_file[15][7]  ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   CLKBUFX2M FE_OFC33_REG0_2_ (.Y(REG0[2]), 
	.A(FE_OFN33_REG0_2_));
   BUFX8M FE_OFC32_REG0_3_ (.Y(REG0[3]), 
	.A(FE_OFN32_REG0_3_));
   BUFX8M FE_OFC31_REG0_4_ (.Y(REG0[4]), 
	.A(FE_OFN31_REG0_4_));
   BUFX10M FE_OFC30_REG0_5_ (.Y(REG0[5]), 
	.A(FE_OFN30_REG0_5_));
   BUFX10M FE_OFC29_REG0_6_ (.Y(REG0[6]), 
	.A(FE_OFN29_REG0_6_));
   BUFX10M FE_OFC28_REG0_7_ (.Y(REG0[7]), 
	.A(FE_OFN28_REG0_7_));
   BUFX8M FE_OFC27_REG1_7_ (.Y(REG1[7]), 
	.A(FE_OFN27_REG1_7_));
   BUFX8M FE_OFC26_REG1_6_ (.Y(REG1[6]), 
	.A(FE_OFN26_REG1_6_));
   BUFX4M FE_OFC25_SE (.Y(FE_OFN25_SE), 
	.A(FE_OFN19_SE));
   SDFFRQX2M \reg_file_reg[5][7]  (.SI(\reg_file[5][6] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[5][7] ), 
	.D(n248), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[5][6]  (.SI(\reg_file[5][5] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[5][6] ), 
	.D(n247), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[5][5]  (.SI(\reg_file[5][4] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[5][5] ), 
	.D(n246), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[5][4]  (.SI(\reg_file[5][3] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[5][4] ), 
	.D(n245), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[5][3]  (.SI(\reg_file[5][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[5][3] ), 
	.D(n244), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[5][2]  (.SI(\reg_file[5][1] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[5][2] ), 
	.D(n243), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[5][1]  (.SI(\reg_file[5][0] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[5][1] ), 
	.D(n242), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[5][0]  (.SI(\reg_file[4][7] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[5][0] ), 
	.D(n241), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[9][7]  (.SI(\reg_file[9][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[9][7] ), 
	.D(n216), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[9][6]  (.SI(\reg_file[9][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[9][6] ), 
	.D(n215), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[9][5]  (.SI(\reg_file[9][4] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[9][5] ), 
	.D(n214), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[9][4]  (.SI(\reg_file[9][3] ), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[9][4] ), 
	.D(n213), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[9][3]  (.SI(\reg_file[9][2] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\reg_file[9][3] ), 
	.D(n212), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[9][2]  (.SI(\reg_file[9][1] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[9][2] ), 
	.D(n211), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[9][1]  (.SI(\reg_file[9][0] ), 
	.SE(FE_OFN19_SE), 
	.RN(RST_n), 
	.Q(\reg_file[9][1] ), 
	.D(n210), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[9][0]  (.SI(\reg_file[8][7] ), 
	.SE(FE_OFN22_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[9][0] ), 
	.D(n209), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[13][7]  (.SI(\reg_file[13][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[13][7] ), 
	.D(n184), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[13][6]  (.SI(\reg_file[13][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[13][6] ), 
	.D(n183), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[13][5]  (.SI(\reg_file[13][4] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[13][5] ), 
	.D(n182), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[13][4]  (.SI(\reg_file[13][3] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[13][4] ), 
	.D(n181), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[13][3]  (.SI(\reg_file[13][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[13][3] ), 
	.D(n180), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[13][2]  (.SI(\reg_file[13][1] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[13][2] ), 
	.D(n179), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[13][1]  (.SI(\reg_file[13][0] ), 
	.SE(FE_OFN22_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[13][1] ), 
	.D(n178), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[13][0]  (.SI(\reg_file[12][7] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[13][0] ), 
	.D(n177), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[7][7]  (.SI(\reg_file[7][6] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[7][7] ), 
	.D(n232), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[7][6]  (.SI(\reg_file[7][5] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[7][6] ), 
	.D(n231), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[7][5]  (.SI(\reg_file[7][4] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[7][5] ), 
	.D(n230), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[7][4]  (.SI(\reg_file[7][3] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[7][4] ), 
	.D(n229), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[7][3]  (.SI(\reg_file[7][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[7][3] ), 
	.D(n228), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[7][2]  (.SI(\reg_file[7][1] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[7][2] ), 
	.D(n227), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[7][1]  (.SI(\reg_file[7][0] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[7][1] ), 
	.D(n226), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[7][0]  (.SI(\reg_file[6][7] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[7][0] ), 
	.D(n225), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[11][7]  (.SI(\reg_file[11][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[11][7] ), 
	.D(n200), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[11][6]  (.SI(\reg_file[11][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[11][6] ), 
	.D(n199), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[11][5]  (.SI(test_si2), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[11][5] ), 
	.D(n198), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[11][4]  (.SI(\reg_file[11][3] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[11][4] ), 
	.D(n197), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[11][3]  (.SI(\reg_file[11][2] ), 
	.SE(FE_OFN19_SE), 
	.RN(RST_n), 
	.Q(\reg_file[11][3] ), 
	.D(n196), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[11][2]  (.SI(\reg_file[11][1] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[11][2] ), 
	.D(n195), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[11][1]  (.SI(\reg_file[11][0] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[11][1] ), 
	.D(n194), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[11][0]  (.SI(\reg_file[10][7] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[11][0] ), 
	.D(n193), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[15][7]  (.SI(\reg_file[15][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[15][7] ), 
	.D(n168), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[15][6]  (.SI(\reg_file[15][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[15][6] ), 
	.D(n167), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[15][5]  (.SI(\reg_file[15][4] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[15][5] ), 
	.D(n166), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[15][4]  (.SI(\reg_file[15][3] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[15][4] ), 
	.D(n165), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[15][3]  (.SI(\reg_file[15][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[15][3] ), 
	.D(n164), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[15][2]  (.SI(\reg_file[15][1] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[15][2] ), 
	.D(n163), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[15][1]  (.SI(\reg_file[15][0] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[15][1] ), 
	.D(n162), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[15][0]  (.SI(\reg_file[14][7] ), 
	.SE(FE_OFN22_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[15][0] ), 
	.D(n161), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[6][7]  (.SI(\reg_file[6][6] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[6][7] ), 
	.D(n240), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[6][6]  (.SI(\reg_file[6][5] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[6][6] ), 
	.D(n239), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[6][5]  (.SI(\reg_file[6][4] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[6][5] ), 
	.D(n238), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[6][4]  (.SI(\reg_file[6][3] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[6][4] ), 
	.D(n237), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[6][3]  (.SI(\reg_file[6][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[6][3] ), 
	.D(n236), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[6][2]  (.SI(\reg_file[6][1] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[6][2] ), 
	.D(n235), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[6][1]  (.SI(\reg_file[6][0] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[6][1] ), 
	.D(n234), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[6][0]  (.SI(\reg_file[5][7] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[6][0] ), 
	.D(n233), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[10][7]  (.SI(\reg_file[10][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[10][7] ), 
	.D(n208), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[10][6]  (.SI(\reg_file[10][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[10][6] ), 
	.D(n207), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[10][5]  (.SI(\reg_file[10][4] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[10][5] ), 
	.D(n206), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[10][4]  (.SI(\reg_file[10][3] ), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[10][4] ), 
	.D(n205), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[10][3]  (.SI(\reg_file[10][2] ), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[10][3] ), 
	.D(n204), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[10][2]  (.SI(\reg_file[10][1] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[10][2] ), 
	.D(n203), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[10][1]  (.SI(\reg_file[10][0] ), 
	.SE(FE_OFN19_SE), 
	.RN(RST_n), 
	.Q(\reg_file[10][1] ), 
	.D(n202), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[10][0]  (.SI(\reg_file[9][7] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[10][0] ), 
	.D(n201), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[14][7]  (.SI(\reg_file[14][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[14][7] ), 
	.D(n176), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[14][6]  (.SI(\reg_file[14][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[14][6] ), 
	.D(n175), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[14][5]  (.SI(\reg_file[14][4] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[14][5] ), 
	.D(n174), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[14][4]  (.SI(\reg_file[14][3] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[14][4] ), 
	.D(n173), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[14][3]  (.SI(\reg_file[14][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[14][3] ), 
	.D(n172), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[14][2]  (.SI(\reg_file[14][1] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[14][2] ), 
	.D(n171), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[14][1]  (.SI(\reg_file[14][0] ), 
	.SE(FE_OFN22_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[14][1] ), 
	.D(n170), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[14][0]  (.SI(\reg_file[13][7] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[14][0] ), 
	.D(n169), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[4][7]  (.SI(\reg_file[4][6] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[4][7] ), 
	.D(n256), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[4][6]  (.SI(\reg_file[4][5] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[4][6] ), 
	.D(n255), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[4][5]  (.SI(\reg_file[4][4] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN10_RST_D1_M), 
	.Q(\reg_file[4][5] ), 
	.D(n254), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[4][4]  (.SI(\reg_file[4][3] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[4][4] ), 
	.D(n253), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[4][3]  (.SI(\reg_file[4][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[4][3] ), 
	.D(n252), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[4][2]  (.SI(\reg_file[4][1] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[4][2] ), 
	.D(n251), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[4][1]  (.SI(\reg_file[4][0] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[4][1] ), 
	.D(n250), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[4][0]  (.SI(REG1[7]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\reg_file[4][0] ), 
	.D(n249), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[8][7]  (.SI(\reg_file[8][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[8][7] ), 
	.D(n224), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[8][6]  (.SI(\reg_file[8][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[8][6] ), 
	.D(n223), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[8][5]  (.SI(\reg_file[8][4] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[8][5] ), 
	.D(n222), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[8][4]  (.SI(\reg_file[8][3] ), 
	.SE(FE_OFN19_SE), 
	.RN(RST_n), 
	.Q(\reg_file[8][4] ), 
	.D(n221), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[8][3]  (.SI(\reg_file[8][2] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[8][3] ), 
	.D(n220), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \reg_file_reg[8][2]  (.SI(\reg_file[8][1] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[8][2] ), 
	.D(n219), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \reg_file_reg[8][1]  (.SI(\reg_file[8][0] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[8][1] ), 
	.D(n218), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[8][0]  (.SI(\reg_file[7][7] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[8][0] ), 
	.D(n217), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[12][7]  (.SI(\reg_file[12][6] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[12][7] ), 
	.D(n192), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[12][6]  (.SI(\reg_file[12][5] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[12][6] ), 
	.D(n191), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[12][5]  (.SI(\reg_file[12][4] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[12][5] ), 
	.D(n190), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[12][4]  (.SI(\reg_file[12][3] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[12][4] ), 
	.D(n189), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[12][3]  (.SI(\reg_file[12][2] ), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[12][3] ), 
	.D(n188), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[12][2]  (.SI(\reg_file[12][1] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[12][2] ), 
	.D(n187), 
	.CK(REF_CLK_M__L5_N5));
   SDFFRQX2M \reg_file_reg[12][1]  (.SI(\reg_file[12][0] ), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(\reg_file[12][1] ), 
	.D(n186), 
	.CK(CLK));
   SDFFRQX2M \reg_file_reg[12][0]  (.SI(\reg_file[11][7] ), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(\reg_file[12][0] ), 
	.D(n185), 
	.CK(CLK));
   SDFFRQX2M \RdData_reg[7]  (.SI(RdData[6]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(RdData[7]), 
	.D(n280), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \RdData_reg[6]  (.SI(RdData[5]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(RdData[6]), 
	.D(n279), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \RdData_reg[5]  (.SI(RdData[4]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(RdData[5]), 
	.D(n278), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \RdData_reg[4]  (.SI(RdData[3]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(RdData[4]), 
	.D(n277), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \RdData_reg[3]  (.SI(RdData[2]), 
	.SE(test_se), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(RdData[3]), 
	.D(n276), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \RdData_reg[2]  (.SI(RdData[1]), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(RdData[2]), 
	.D(n275), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \RdData_reg[1]  (.SI(RdData[0]), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(RdData[1]), 
	.D(n274), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \RdData_reg[0]  (.SI(RdData_Valid), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(RdData[0]), 
	.D(n273), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M RdData_Valid_reg (.SI(test_si1), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(RdData_Valid), 
	.D(n376), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \reg_file_reg[0][0]  (.SI(RdData[7]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(REG0[0]), 
	.D(n265), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \reg_file_reg[0][1]  (.SI(n348), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(REG0[1]), 
	.D(n266), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRQX2M \reg_file_reg[0][2]  (.SI(REG0[1]), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(FE_OFN33_REG0_2_), 
	.D(n267), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX2M \reg_file_reg[0][3]  (.SI(REG0[2]), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(FE_OFN32_REG0_3_), 
	.D(n268), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX2M \reg_file_reg[0][4]  (.SI(REG0[3]), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(FE_OFN31_REG0_4_), 
	.D(n269), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX2M \reg_file_reg[0][5]  (.SI(REG0[4]), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(FE_OFN30_REG0_5_), 
	.D(n270), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX2M \reg_file_reg[0][6]  (.SI(REG0[5]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN8_RST_D1_M), 
	.Q(FE_OFN29_REG0_6_), 
	.D(n271), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRHQX2M \reg_file_reg[0][7]  (.SI(n349), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(FE_OFN28_REG0_7_), 
	.D(n272), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX4M \reg_file_reg[1][5]  (.SI(REG1[4]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(REG1[5]), 
	.D(n262), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRHQX4M \reg_file_reg[1][4]  (.SI(REG1[3]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(REG1[4]), 
	.D(n261), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX4M \reg_file_reg[1][1]  (.SI(REG1[0]), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(REG1[1]), 
	.D(n258), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX2M \reg_file_reg[1][7]  (.SI(REG1[6]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(FE_OFN27_REG1_7_), 
	.D(n264), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRHQX4M \reg_file_reg[1][3]  (.SI(REG1[2]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(REG1[3]), 
	.D(n260), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX4M \reg_file_reg[1][2]  (.SI(REG1[1]), 
	.SE(FE_OFN25_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(REG1[2]), 
	.D(n259), 
	.CK(REF_CLK_M__L5_N6));
   SDFFRHQX2M \reg_file_reg[1][6]  (.SI(n347), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(FE_OFN26_REG1_6_), 
	.D(n263), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRHQX4M \reg_file_reg[1][0]  (.SI(REG0[7]), 
	.SE(FE_OFN19_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(REG1[0]), 
	.D(n257), 
	.CK(REF_CLK_M__L5_N6));
   AND2X2M U172 (.Y(n299), 
	.B(REG1[0]), 
	.A(N10));
   AND2X2M U173 (.Y(n300), 
	.B(REG1[6]), 
	.A(N10));
   INVX6M U174 (.Y(n357), 
	.A(n358));
   NAND2X2M U182 (.Y(n146), 
	.B(n138), 
	.A(n147));
   NAND2X2M U183 (.Y(n148), 
	.B(n140), 
	.A(n147));
   NAND2X2M U184 (.Y(n149), 
	.B(n142), 
	.A(n147));
   NAND2X2M U185 (.Y(n150), 
	.B(n144), 
	.A(n147));
   NAND2X2M U186 (.Y(n157), 
	.B(n357), 
	.A(n158));
   NOR2X2M U187 (.Y(n144), 
	.B(N11), 
	.A(n357));
   AOI31X2M U198 (.Y(n151), 
	.B0(n379), 
	.A2(n377), 
	.A1(n378), 
	.A0(N11));
   NAND2X2M U199 (.Y(n139), 
	.B(n137), 
	.A(n140));
   NAND2X2M U200 (.Y(n141), 
	.B(n137), 
	.A(n142));
   NAND2X2M U201 (.Y(n143), 
	.B(n137), 
	.A(n144));
   NAND2X2M U202 (.Y(n152), 
	.B(n138), 
	.A(n153));
   NAND2X2M U203 (.Y(n154), 
	.B(n140), 
	.A(n153));
   NAND2X2M U204 (.Y(n155), 
	.B(n142), 
	.A(n153));
   NAND2X2M U205 (.Y(n156), 
	.B(n144), 
	.A(n153));
   NAND2X2M U206 (.Y(n159), 
	.B(n358), 
	.A(n158));
   NAND2X2M U207 (.Y(n136), 
	.B(n138), 
	.A(n137));
   AND3X2M U208 (.Y(n158), 
	.C(n378), 
	.B(n377), 
	.A(n151));
   AND2X2M U209 (.Y(n147), 
	.B(n377), 
	.A(n145));
   NOR2X2M U210 (.Y(n138), 
	.B(n359), 
	.A(n358));
   NOR2X2M U211 (.Y(n142), 
	.B(N11), 
	.A(n358));
   NOR2X2M U212 (.Y(n140), 
	.B(n357), 
	.A(n359));
   INVX2M U213 (.Y(n380), 
	.A(WrData[0]));
   INVX2M U214 (.Y(n381), 
	.A(WrData[1]));
   INVX2M U215 (.Y(n382), 
	.A(WrData[2]));
   INVX2M U216 (.Y(n383), 
	.A(WrData[3]));
   INVX2M U217 (.Y(n384), 
	.A(WrData[4]));
   INVX2M U218 (.Y(n385), 
	.A(WrData[5]));
   INVX2M U219 (.Y(n386), 
	.A(WrData[6]));
   INVX2M U220 (.Y(n376), 
	.A(n160));
   AND3X2M U225 (.Y(n153), 
	.C(N12), 
	.B(n378), 
	.A(n151));
   INVX2M U226 (.Y(n378), 
	.A(N13));
   AND2X2M U227 (.Y(n137), 
	.B(N12), 
	.A(n145));
   INVX2M U228 (.Y(n377), 
	.A(N12));
   AND2X2M U229 (.Y(n145), 
	.B(N13), 
	.A(n151));
   INVX2M U230 (.Y(n358), 
	.A(N10));
   INVX2M U231 (.Y(n359), 
	.A(N11));
   INVX2M U232 (.Y(n387), 
	.A(WrData[7]));
   NAND2X2M U233 (.Y(n160), 
	.B(n379), 
	.A(RdEn));
   INVX2M U234 (.Y(n379), 
	.A(WrEn));
   MXI2X1M U237 (.Y(n346), 
	.S0(N11), 
	.B(N10), 
	.A(n345));
   NOR2BX2M U238 (.Y(n345), 
	.B(N10), 
	.AN(REG0[5]));
   MXI2X1M U239 (.Y(n344), 
	.S0(N11), 
	.B(n358), 
	.A(n299));
   MXI2X1M U240 (.Y(n335), 
	.S0(N11), 
	.B(n358), 
	.A(n300));
   OAI2BB2X1M U241 (.Y(n225), 
	.B1(n152), 
	.B0(n380), 
	.A1N(n152), 
	.A0N(\reg_file[7][0] ));
   OAI2BB2X1M U242 (.Y(n226), 
	.B1(n152), 
	.B0(n381), 
	.A1N(n152), 
	.A0N(\reg_file[7][1] ));
   OAI2BB2X1M U243 (.Y(n227), 
	.B1(n152), 
	.B0(n382), 
	.A1N(n152), 
	.A0N(\reg_file[7][2] ));
   OAI2BB2X1M U244 (.Y(n228), 
	.B1(n152), 
	.B0(n383), 
	.A1N(n152), 
	.A0N(\reg_file[7][3] ));
   OAI2BB2X1M U245 (.Y(n229), 
	.B1(n152), 
	.B0(n384), 
	.A1N(n152), 
	.A0N(\reg_file[7][4] ));
   OAI2BB2X1M U246 (.Y(n230), 
	.B1(n152), 
	.B0(n385), 
	.A1N(n152), 
	.A0N(\reg_file[7][5] ));
   OAI2BB2X1M U247 (.Y(n231), 
	.B1(n152), 
	.B0(n386), 
	.A1N(n152), 
	.A0N(\reg_file[7][6] ));
   OAI2BB2X1M U248 (.Y(n232), 
	.B1(n152), 
	.B0(n387), 
	.A1N(n152), 
	.A0N(\reg_file[7][7] ));
   OAI2BB2X1M U249 (.Y(n233), 
	.B1(n154), 
	.B0(n380), 
	.A1N(n154), 
	.A0N(\reg_file[6][0] ));
   OAI2BB2X1M U250 (.Y(n234), 
	.B1(n154), 
	.B0(n381), 
	.A1N(n154), 
	.A0N(\reg_file[6][1] ));
   OAI2BB2X1M U251 (.Y(n235), 
	.B1(n154), 
	.B0(n382), 
	.A1N(n154), 
	.A0N(\reg_file[6][2] ));
   OAI2BB2X1M U252 (.Y(n236), 
	.B1(n154), 
	.B0(n383), 
	.A1N(n154), 
	.A0N(\reg_file[6][3] ));
   OAI2BB2X1M U253 (.Y(n237), 
	.B1(n154), 
	.B0(n384), 
	.A1N(n154), 
	.A0N(\reg_file[6][4] ));
   OAI2BB2X1M U254 (.Y(n238), 
	.B1(n154), 
	.B0(n385), 
	.A1N(n154), 
	.A0N(\reg_file[6][5] ));
   OAI2BB2X1M U255 (.Y(n239), 
	.B1(n154), 
	.B0(n386), 
	.A1N(n154), 
	.A0N(\reg_file[6][6] ));
   OAI2BB2X1M U256 (.Y(n240), 
	.B1(n154), 
	.B0(n387), 
	.A1N(n154), 
	.A0N(\reg_file[6][7] ));
   OAI2BB2X1M U257 (.Y(n241), 
	.B1(n155), 
	.B0(n380), 
	.A1N(n155), 
	.A0N(\reg_file[5][0] ));
   OAI2BB2X1M U258 (.Y(n242), 
	.B1(n155), 
	.B0(n381), 
	.A1N(n155), 
	.A0N(\reg_file[5][1] ));
   OAI2BB2X1M U259 (.Y(n243), 
	.B1(n155), 
	.B0(n382), 
	.A1N(n155), 
	.A0N(\reg_file[5][2] ));
   OAI2BB2X1M U260 (.Y(n244), 
	.B1(n155), 
	.B0(n383), 
	.A1N(n155), 
	.A0N(\reg_file[5][3] ));
   OAI2BB2X1M U261 (.Y(n245), 
	.B1(n155), 
	.B0(n384), 
	.A1N(n155), 
	.A0N(\reg_file[5][4] ));
   OAI2BB2X1M U262 (.Y(n246), 
	.B1(n155), 
	.B0(n385), 
	.A1N(n155), 
	.A0N(\reg_file[5][5] ));
   OAI2BB2X1M U263 (.Y(n247), 
	.B1(n155), 
	.B0(n386), 
	.A1N(n155), 
	.A0N(\reg_file[5][6] ));
   OAI2BB2X1M U264 (.Y(n248), 
	.B1(n155), 
	.B0(n387), 
	.A1N(n155), 
	.A0N(\reg_file[5][7] ));
   OAI2BB2X1M U265 (.Y(n249), 
	.B1(n156), 
	.B0(n380), 
	.A1N(n156), 
	.A0N(\reg_file[4][0] ));
   OAI2BB2X1M U266 (.Y(n250), 
	.B1(n156), 
	.B0(n381), 
	.A1N(n156), 
	.A0N(\reg_file[4][1] ));
   OAI2BB2X1M U267 (.Y(n251), 
	.B1(n156), 
	.B0(n382), 
	.A1N(n156), 
	.A0N(\reg_file[4][2] ));
   OAI2BB2X1M U268 (.Y(n252), 
	.B1(n156), 
	.B0(n383), 
	.A1N(n156), 
	.A0N(\reg_file[4][3] ));
   OAI2BB2X1M U269 (.Y(n253), 
	.B1(n156), 
	.B0(n384), 
	.A1N(n156), 
	.A0N(\reg_file[4][4] ));
   OAI2BB2X1M U270 (.Y(n254), 
	.B1(n156), 
	.B0(n385), 
	.A1N(n156), 
	.A0N(\reg_file[4][5] ));
   OAI2BB2X1M U271 (.Y(n255), 
	.B1(n156), 
	.B0(n386), 
	.A1N(n156), 
	.A0N(\reg_file[4][6] ));
   OAI2BB2X1M U272 (.Y(n256), 
	.B1(n156), 
	.B0(n387), 
	.A1N(n156), 
	.A0N(\reg_file[4][7] ));
   OAI2BB2X1M U273 (.Y(n169), 
	.B1(n139), 
	.B0(n380), 
	.A1N(n139), 
	.A0N(\reg_file[14][0] ));
   OAI2BB2X1M U274 (.Y(n170), 
	.B1(n139), 
	.B0(n381), 
	.A1N(n139), 
	.A0N(\reg_file[14][1] ));
   OAI2BB2X1M U275 (.Y(n171), 
	.B1(n139), 
	.B0(n382), 
	.A1N(n139), 
	.A0N(\reg_file[14][2] ));
   OAI2BB2X1M U276 (.Y(n172), 
	.B1(n139), 
	.B0(n383), 
	.A1N(n139), 
	.A0N(\reg_file[14][3] ));
   OAI2BB2X1M U277 (.Y(n173), 
	.B1(n139), 
	.B0(n384), 
	.A1N(n139), 
	.A0N(\reg_file[14][4] ));
   OAI2BB2X1M U278 (.Y(n174), 
	.B1(n139), 
	.B0(n385), 
	.A1N(n139), 
	.A0N(\reg_file[14][5] ));
   OAI2BB2X1M U279 (.Y(n175), 
	.B1(n139), 
	.B0(n386), 
	.A1N(n139), 
	.A0N(\reg_file[14][6] ));
   OAI2BB2X1M U280 (.Y(n176), 
	.B1(n139), 
	.B0(n387), 
	.A1N(n139), 
	.A0N(\reg_file[14][7] ));
   OAI2BB2X1M U281 (.Y(n177), 
	.B1(n141), 
	.B0(n380), 
	.A1N(n141), 
	.A0N(\reg_file[13][0] ));
   OAI2BB2X1M U282 (.Y(n178), 
	.B1(n141), 
	.B0(n381), 
	.A1N(n141), 
	.A0N(\reg_file[13][1] ));
   OAI2BB2X1M U283 (.Y(n179), 
	.B1(n141), 
	.B0(n382), 
	.A1N(n141), 
	.A0N(\reg_file[13][2] ));
   OAI2BB2X1M U284 (.Y(n180), 
	.B1(n141), 
	.B0(n383), 
	.A1N(n141), 
	.A0N(\reg_file[13][3] ));
   OAI2BB2X1M U285 (.Y(n181), 
	.B1(n141), 
	.B0(n384), 
	.A1N(n141), 
	.A0N(\reg_file[13][4] ));
   OAI2BB2X1M U286 (.Y(n182), 
	.B1(n141), 
	.B0(n385), 
	.A1N(n141), 
	.A0N(\reg_file[13][5] ));
   OAI2BB2X1M U287 (.Y(n183), 
	.B1(n141), 
	.B0(n386), 
	.A1N(n141), 
	.A0N(\reg_file[13][6] ));
   OAI2BB2X1M U288 (.Y(n184), 
	.B1(n141), 
	.B0(n387), 
	.A1N(n141), 
	.A0N(\reg_file[13][7] ));
   OAI2BB2X1M U289 (.Y(n185), 
	.B1(n143), 
	.B0(n380), 
	.A1N(n143), 
	.A0N(\reg_file[12][0] ));
   OAI2BB2X1M U290 (.Y(n186), 
	.B1(n143), 
	.B0(n381), 
	.A1N(n143), 
	.A0N(\reg_file[12][1] ));
   OAI2BB2X1M U291 (.Y(n187), 
	.B1(n143), 
	.B0(n382), 
	.A1N(n143), 
	.A0N(\reg_file[12][2] ));
   OAI2BB2X1M U292 (.Y(n188), 
	.B1(n143), 
	.B0(n383), 
	.A1N(n143), 
	.A0N(\reg_file[12][3] ));
   OAI2BB2X1M U293 (.Y(n189), 
	.B1(n143), 
	.B0(n384), 
	.A1N(n143), 
	.A0N(\reg_file[12][4] ));
   OAI2BB2X1M U294 (.Y(n190), 
	.B1(n143), 
	.B0(n385), 
	.A1N(n143), 
	.A0N(\reg_file[12][5] ));
   OAI2BB2X1M U295 (.Y(n191), 
	.B1(n143), 
	.B0(n386), 
	.A1N(n143), 
	.A0N(\reg_file[12][6] ));
   OAI2BB2X1M U296 (.Y(n192), 
	.B1(n143), 
	.B0(n387), 
	.A1N(n143), 
	.A0N(\reg_file[12][7] ));
   OAI2BB2X1M U297 (.Y(n161), 
	.B1(n380), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][0] ));
   OAI2BB2X1M U298 (.Y(n162), 
	.B1(n381), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][1] ));
   OAI2BB2X1M U299 (.Y(n163), 
	.B1(n382), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][2] ));
   OAI2BB2X1M U300 (.Y(n164), 
	.B1(n383), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][3] ));
   OAI2BB2X1M U301 (.Y(n165), 
	.B1(n384), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][4] ));
   OAI2BB2X1M U302 (.Y(n166), 
	.B1(n385), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][5] ));
   OAI2BB2X1M U303 (.Y(n167), 
	.B1(n386), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][6] ));
   OAI2BB2X1M U304 (.Y(n168), 
	.B1(n387), 
	.B0(n136), 
	.A1N(n136), 
	.A0N(\reg_file[15][7] ));
   OAI2BB2X1M U305 (.Y(n193), 
	.B1(n146), 
	.B0(n380), 
	.A1N(n146), 
	.A0N(\reg_file[11][0] ));
   OAI2BB2X1M U306 (.Y(n194), 
	.B1(n146), 
	.B0(n381), 
	.A1N(n146), 
	.A0N(\reg_file[11][1] ));
   OAI2BB2X1M U307 (.Y(n195), 
	.B1(n146), 
	.B0(n382), 
	.A1N(n146), 
	.A0N(\reg_file[11][2] ));
   OAI2BB2X1M U308 (.Y(n196), 
	.B1(n146), 
	.B0(n383), 
	.A1N(n146), 
	.A0N(\reg_file[11][3] ));
   OAI2BB2X1M U309 (.Y(n197), 
	.B1(n146), 
	.B0(n384), 
	.A1N(n146), 
	.A0N(\reg_file[11][4] ));
   OAI2BB2X1M U310 (.Y(n198), 
	.B1(n146), 
	.B0(n385), 
	.A1N(n146), 
	.A0N(\reg_file[11][5] ));
   OAI2BB2X1M U311 (.Y(n199), 
	.B1(n146), 
	.B0(n386), 
	.A1N(n146), 
	.A0N(\reg_file[11][6] ));
   OAI2BB2X1M U312 (.Y(n200), 
	.B1(n146), 
	.B0(n387), 
	.A1N(n146), 
	.A0N(\reg_file[11][7] ));
   OAI2BB2X1M U313 (.Y(n201), 
	.B1(n148), 
	.B0(n380), 
	.A1N(n148), 
	.A0N(\reg_file[10][0] ));
   OAI2BB2X1M U314 (.Y(n202), 
	.B1(n148), 
	.B0(n381), 
	.A1N(n148), 
	.A0N(\reg_file[10][1] ));
   OAI2BB2X1M U315 (.Y(n203), 
	.B1(n148), 
	.B0(n382), 
	.A1N(n148), 
	.A0N(\reg_file[10][2] ));
   OAI2BB2X1M U316 (.Y(n204), 
	.B1(n148), 
	.B0(n383), 
	.A1N(n148), 
	.A0N(\reg_file[10][3] ));
   OAI2BB2X1M U317 (.Y(n205), 
	.B1(n148), 
	.B0(n384), 
	.A1N(n148), 
	.A0N(\reg_file[10][4] ));
   OAI2BB2X1M U318 (.Y(n206), 
	.B1(n148), 
	.B0(n385), 
	.A1N(n148), 
	.A0N(\reg_file[10][5] ));
   OAI2BB2X1M U319 (.Y(n207), 
	.B1(n148), 
	.B0(n386), 
	.A1N(n148), 
	.A0N(\reg_file[10][6] ));
   OAI2BB2X1M U320 (.Y(n208), 
	.B1(n148), 
	.B0(n387), 
	.A1N(n148), 
	.A0N(\reg_file[10][7] ));
   OAI2BB2X1M U321 (.Y(n209), 
	.B1(n149), 
	.B0(n380), 
	.A1N(n149), 
	.A0N(\reg_file[9][0] ));
   OAI2BB2X1M U322 (.Y(n210), 
	.B1(n149), 
	.B0(n381), 
	.A1N(n149), 
	.A0N(\reg_file[9][1] ));
   OAI2BB2X1M U323 (.Y(n211), 
	.B1(n149), 
	.B0(n382), 
	.A1N(n149), 
	.A0N(\reg_file[9][2] ));
   OAI2BB2X1M U324 (.Y(n212), 
	.B1(n149), 
	.B0(n383), 
	.A1N(n149), 
	.A0N(\reg_file[9][3] ));
   OAI2BB2X1M U325 (.Y(n213), 
	.B1(n149), 
	.B0(n384), 
	.A1N(n149), 
	.A0N(\reg_file[9][4] ));
   OAI2BB2X1M U326 (.Y(n214), 
	.B1(n149), 
	.B0(n385), 
	.A1N(n149), 
	.A0N(\reg_file[9][5] ));
   OAI2BB2X1M U327 (.Y(n215), 
	.B1(n149), 
	.B0(n386), 
	.A1N(n149), 
	.A0N(\reg_file[9][6] ));
   OAI2BB2X1M U328 (.Y(n216), 
	.B1(n149), 
	.B0(n387), 
	.A1N(n149), 
	.A0N(\reg_file[9][7] ));
   OAI2BB2X1M U329 (.Y(n217), 
	.B1(n150), 
	.B0(n380), 
	.A1N(n150), 
	.A0N(\reg_file[8][0] ));
   OAI2BB2X1M U330 (.Y(n218), 
	.B1(n150), 
	.B0(n381), 
	.A1N(n150), 
	.A0N(\reg_file[8][1] ));
   OAI2BB2X1M U331 (.Y(n219), 
	.B1(n150), 
	.B0(n382), 
	.A1N(n150), 
	.A0N(\reg_file[8][2] ));
   OAI2BB2X1M U332 (.Y(n220), 
	.B1(n150), 
	.B0(n383), 
	.A1N(n150), 
	.A0N(\reg_file[8][3] ));
   OAI2BB2X1M U333 (.Y(n221), 
	.B1(n150), 
	.B0(n384), 
	.A1N(n150), 
	.A0N(\reg_file[8][4] ));
   OAI2BB2X1M U334 (.Y(n222), 
	.B1(n150), 
	.B0(n385), 
	.A1N(n150), 
	.A0N(\reg_file[8][5] ));
   OAI2BB2X1M U335 (.Y(n223), 
	.B1(n150), 
	.B0(n386), 
	.A1N(n150), 
	.A0N(\reg_file[8][6] ));
   OAI2BB2X1M U336 (.Y(n224), 
	.B1(n150), 
	.B0(n387), 
	.A1N(n150), 
	.A0N(\reg_file[8][7] ));
   OAI2BB2X1M U337 (.Y(n257), 
	.B1(n157), 
	.B0(n380), 
	.A1N(n157), 
	.A0N(REG1[0]));
   OAI2BB2X1M U338 (.Y(n258), 
	.B1(n157), 
	.B0(n381), 
	.A1N(n157), 
	.A0N(REG1[1]));
   OAI2BB2X1M U339 (.Y(n259), 
	.B1(n157), 
	.B0(n382), 
	.A1N(n157), 
	.A0N(REG1[2]));
   OAI2BB2X1M U340 (.Y(n260), 
	.B1(n157), 
	.B0(n383), 
	.A1N(n157), 
	.A0N(REG1[3]));
   OAI2BB2X1M U341 (.Y(n261), 
	.B1(n157), 
	.B0(n384), 
	.A1N(n157), 
	.A0N(REG1[4]));
   OAI2BB2X1M U342 (.Y(n262), 
	.B1(n157), 
	.B0(n385), 
	.A1N(n157), 
	.A0N(REG1[5]));
   OAI2BB2X1M U343 (.Y(n263), 
	.B1(n157), 
	.B0(n386), 
	.A1N(n157), 
	.A0N(REG1[6]));
   OAI2BB2X1M U344 (.Y(n264), 
	.B1(n157), 
	.B0(n387), 
	.A1N(n157), 
	.A0N(REG1[7]));
   OAI2BB2X1M U345 (.Y(n265), 
	.B1(n159), 
	.B0(n380), 
	.A1N(n159), 
	.A0N(REG0[0]));
   OAI2BB2X1M U346 (.Y(n266), 
	.B1(n159), 
	.B0(n381), 
	.A1N(n159), 
	.A0N(REG0[1]));
   OAI2BB2X1M U347 (.Y(n267), 
	.B1(n159), 
	.B0(n382), 
	.A1N(n159), 
	.A0N(REG0[2]));
   OAI2BB2X1M U348 (.Y(n268), 
	.B1(n159), 
	.B0(n383), 
	.A1N(n159), 
	.A0N(REG0[3]));
   OAI2BB2X1M U349 (.Y(n269), 
	.B1(n159), 
	.B0(n384), 
	.A1N(n159), 
	.A0N(REG0[4]));
   OAI2BB2X1M U350 (.Y(n270), 
	.B1(n159), 
	.B0(n385), 
	.A1N(n159), 
	.A0N(REG0[5]));
   OAI2BB2X1M U351 (.Y(n271), 
	.B1(n159), 
	.B0(n386), 
	.A1N(n159), 
	.A0N(REG0[6]));
   OAI2BB2X1M U352 (.Y(n272), 
	.B1(n159), 
	.B0(n387), 
	.A1N(n159), 
	.A0N(REG0[7]));
   AO22X1M U353 (.Y(n273), 
	.B1(n160), 
	.B0(RdData[0]), 
	.A1(n376), 
	.A0(N58));
   MX4X1M U354 (.Y(N58), 
	.S1(N12), 
	.S0(N13), 
	.D(n301), 
	.C(n303), 
	.B(n302), 
	.A(n304));
   OAI21X2M U355 (.Y(n304), 
	.B0(n344), 
	.A1(n348), 
	.A0(N10));
   MX4X1M U356 (.Y(n301), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][0] ), 
	.C(\reg_file[14][0] ), 
	.B(\reg_file[13][0] ), 
	.A(\reg_file[12][0] ));
   AO22X1M U357 (.Y(n274), 
	.B1(n160), 
	.B0(RdData[1]), 
	.A1(n376), 
	.A0(N57));
   MX4X1M U358 (.Y(N57), 
	.S1(N12), 
	.S0(N13), 
	.D(n305), 
	.C(n307), 
	.B(n306), 
	.A(n308));
   MXI2X1M U359 (.Y(n308), 
	.S0(N10), 
	.B(n342), 
	.A(n343));
   MX4X1M U360 (.Y(n306), 
	.S1(N11), 
	.S0(N10), 
	.D(\reg_file[11][1] ), 
	.C(\reg_file[10][1] ), 
	.B(\reg_file[9][1] ), 
	.A(\reg_file[8][1] ));
   AO22X1M U361 (.Y(n275), 
	.B1(n160), 
	.B0(RdData[2]), 
	.A1(n376), 
	.A0(N56));
   MX4X1M U362 (.Y(N56), 
	.S1(N12), 
	.S0(N13), 
	.D(n309), 
	.C(n311), 
	.B(n310), 
	.A(n312));
   MXI2X1M U363 (.Y(n312), 
	.S0(N10), 
	.B(n340), 
	.A(n341));
   MX4X1M U364 (.Y(n310), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[11][2] ), 
	.C(\reg_file[10][2] ), 
	.B(\reg_file[9][2] ), 
	.A(\reg_file[8][2] ));
   AO22X1M U365 (.Y(n276), 
	.B1(n160), 
	.B0(RdData[3]), 
	.A1(n376), 
	.A0(N55));
   MX4X1M U366 (.Y(N55), 
	.S1(N12), 
	.S0(N13), 
	.D(n313), 
	.C(n315), 
	.B(n314), 
	.A(n316));
   MXI2X1M U367 (.Y(n316), 
	.S0(N10), 
	.B(n338), 
	.A(n339));
   MX4X1M U368 (.Y(n314), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[11][3] ), 
	.C(\reg_file[10][3] ), 
	.B(\reg_file[9][3] ), 
	.A(\reg_file[8][3] ));
   AO22X1M U369 (.Y(n277), 
	.B1(n160), 
	.B0(RdData[4]), 
	.A1(n376), 
	.A0(N54));
   MX4X1M U370 (.Y(N54), 
	.S1(N12), 
	.S0(N13), 
	.D(n317), 
	.C(n319), 
	.B(n318), 
	.A(n320));
   MXI2X1M U371 (.Y(n320), 
	.S0(N10), 
	.B(n336), 
	.A(n337));
   MX4X1M U372 (.Y(n318), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[11][4] ), 
	.C(\reg_file[10][4] ), 
	.B(\reg_file[9][4] ), 
	.A(\reg_file[8][4] ));
   AO22X1M U373 (.Y(n278), 
	.B1(n160), 
	.B0(RdData[5]), 
	.A1(n376), 
	.A0(N53));
   MX4X1M U374 (.Y(N53), 
	.S1(N12), 
	.S0(N13), 
	.D(n321), 
	.C(n323), 
	.B(n322), 
	.A(n324));
   OAI21X2M U375 (.Y(n324), 
	.B0(n346), 
	.A1(n347), 
	.A0(n358));
   MX4X1M U376 (.Y(n322), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[11][5] ), 
	.C(\reg_file[10][5] ), 
	.B(\reg_file[9][5] ), 
	.A(\reg_file[8][5] ));
   AO22X1M U377 (.Y(n279), 
	.B1(n160), 
	.B0(RdData[6]), 
	.A1(n376), 
	.A0(N52));
   MX4X1M U378 (.Y(N52), 
	.S1(N12), 
	.S0(N13), 
	.D(n325), 
	.C(n327), 
	.B(n326), 
	.A(n328));
   OAI21X2M U379 (.Y(n328), 
	.B0(n335), 
	.A1(n349), 
	.A0(N10));
   MX4X1M U380 (.Y(n326), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[11][6] ), 
	.C(\reg_file[10][6] ), 
	.B(\reg_file[9][6] ), 
	.A(\reg_file[8][6] ));
   AO22X1M U381 (.Y(n280), 
	.B1(n160), 
	.B0(RdData[7]), 
	.A1(n376), 
	.A0(N51));
   MX4X1M U382 (.Y(N51), 
	.S1(N12), 
	.S0(N13), 
	.D(n329), 
	.C(n331), 
	.B(n330), 
	.A(n332));
   MXI2X1M U383 (.Y(n332), 
	.S0(N10), 
	.B(n333), 
	.A(n334));
   MX4X1M U384 (.Y(n330), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[11][7] ), 
	.C(\reg_file[10][7] ), 
	.B(\reg_file[9][7] ), 
	.A(\reg_file[8][7] ));
   MX4X1M U385 (.Y(n303), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[7][0] ), 
	.C(\reg_file[6][0] ), 
	.B(\reg_file[5][0] ), 
	.A(\reg_file[4][0] ));
   MX4X1M U386 (.Y(n307), 
	.S1(N11), 
	.S0(N10), 
	.D(\reg_file[7][1] ), 
	.C(\reg_file[6][1] ), 
	.B(\reg_file[5][1] ), 
	.A(\reg_file[4][1] ));
   MX4X1M U387 (.Y(n311), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[7][2] ), 
	.C(\reg_file[6][2] ), 
	.B(\reg_file[5][2] ), 
	.A(\reg_file[4][2] ));
   MX4X1M U388 (.Y(n315), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[7][3] ), 
	.C(\reg_file[6][3] ), 
	.B(\reg_file[5][3] ), 
	.A(\reg_file[4][3] ));
   MX4X1M U389 (.Y(n319), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[7][4] ), 
	.C(\reg_file[6][4] ), 
	.B(\reg_file[5][4] ), 
	.A(\reg_file[4][4] ));
   MX4X1M U390 (.Y(n323), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[7][5] ), 
	.C(\reg_file[6][5] ), 
	.B(\reg_file[5][5] ), 
	.A(\reg_file[4][5] ));
   MX4X1M U391 (.Y(n327), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[7][6] ), 
	.C(\reg_file[6][6] ), 
	.B(\reg_file[5][6] ), 
	.A(\reg_file[4][6] ));
   MX4X1M U392 (.Y(n331), 
	.S1(N11), 
	.S0(N10), 
	.D(\reg_file[7][7] ), 
	.C(\reg_file[6][7] ), 
	.B(\reg_file[5][7] ), 
	.A(\reg_file[4][7] ));
   MX4X1M U393 (.Y(n305), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][1] ), 
	.C(\reg_file[14][1] ), 
	.B(\reg_file[13][1] ), 
	.A(\reg_file[12][1] ));
   MX4X1M U394 (.Y(n309), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][2] ), 
	.C(\reg_file[14][2] ), 
	.B(\reg_file[13][2] ), 
	.A(\reg_file[12][2] ));
   MX4X1M U395 (.Y(n313), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][3] ), 
	.C(\reg_file[14][3] ), 
	.B(\reg_file[13][3] ), 
	.A(\reg_file[12][3] ));
   MX4X1M U396 (.Y(n317), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][4] ), 
	.C(\reg_file[14][4] ), 
	.B(\reg_file[13][4] ), 
	.A(\reg_file[12][4] ));
   MX4X1M U397 (.Y(n321), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][5] ), 
	.C(\reg_file[14][5] ), 
	.B(\reg_file[13][5] ), 
	.A(\reg_file[12][5] ));
   MX4X1M U398 (.Y(n325), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][6] ), 
	.C(\reg_file[14][6] ), 
	.B(\reg_file[13][6] ), 
	.A(\reg_file[12][6] ));
   MX4X1M U399 (.Y(n329), 
	.S1(N11), 
	.S0(n357), 
	.D(\reg_file[15][7] ), 
	.C(\reg_file[14][7] ), 
	.B(\reg_file[13][7] ), 
	.A(\reg_file[12][7] ));
   MX4X1M U400 (.Y(n302), 
	.S1(N11), 
	.S0(N10), 
	.D(\reg_file[11][0] ), 
	.C(\reg_file[10][0] ), 
	.B(\reg_file[9][0] ), 
	.A(\reg_file[8][0] ));
   NAND2X2M U401 (.Y(n340), 
	.B(n359), 
	.A(REG1[2]));
   NAND2X2M U402 (.Y(n338), 
	.B(n359), 
	.A(REG1[3]));
   NAND2X2M U403 (.Y(n333), 
	.B(n359), 
	.A(REG1[7]));
   NAND2X2M U404 (.Y(n342), 
	.B(n359), 
	.A(REG1[1]));
   NAND2X2M U405 (.Y(n336), 
	.B(n359), 
	.A(REG1[4]));
   NAND2X2M U406 (.Y(n343), 
	.B(n359), 
	.A(REG0[1]));
   NAND2X2M U407 (.Y(n341), 
	.B(n359), 
	.A(REG0[2]));
   NAND2X2M U408 (.Y(n339), 
	.B(n359), 
	.A(REG0[3]));
   NAND2X2M U409 (.Y(n337), 
	.B(n359), 
	.A(REG0[4]));
   NAND2X2M U410 (.Y(n334), 
	.B(n359), 
	.A(REG0[7]));
   INVX2M U411 (.Y(n347), 
	.A(REG1[5]));
   INVX2M U412 (.Y(n348), 
	.A(REG0[0]));
   INVX2M U413 (.Y(n349), 
	.A(REG0[6]));
   INVX2M U3 (.Y(REG3[0]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U5 (.Y(REG3[1]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U7 (.Y(REG3[2]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U9 (.Y(REG3[3]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U11 (.Y(REG3[4]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U13 (.Y(REG3[5]), 
	.A(LTIE_LTIELO_NET));
   INVX2M U15 (.Y(REG3[6]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U17 (.Y(REG3[7]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U19 (.Y(REG2[0]), 
	.A(LTIE_LTIELO_NET));
   INVX2M U21 (.Y(REG2[1]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U23 (.Y(REG2[2]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U25 (.Y(REG2[3]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U27 (.Y(REG2[4]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U29 (.Y(REG2[5]), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U31 (.Y(REG2[6]), 
	.A(LTIE_LTIELO_NET));
   INVX2M U33 (.Y(REG2[7]), 
	.A(HTIE_LTIEHI_NET));
endmodule

module ALU_00000008_00000004_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n173, 
	n175, 
	n195);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n173;
   input n175;
   input n195;

   // Internal wires
   wire FE_RN_543_0;
   wire FE_RN_542_0;
   wire FE_RN_541_0;
   wire FE_RN_540_0;
   wire FE_RN_539_0;
   wire FE_RN_538_0;
   wire FE_RN_537_0;
   wire FE_RN_536_0;
   wire FE_RN_535_0;
   wire FE_RN_534_0;
   wire FE_RN_533_0;
   wire FE_RN_532_0;
   wire FE_RN_531_0;
   wire FE_RN_530_0;
   wire FE_RN_529_0;
   wire FE_RN_528_0;
   wire FE_RN_527_0;
   wire FE_RN_526_0;
   wire FE_RN_525_0;
   wire FE_RN_524_0;
   wire FE_RN_523_0;
   wire FE_RN_522_0;
   wire FE_RN_521_0;
   wire FE_RN_520_0;
   wire FE_RN_519_0;
   wire FE_RN_518_0;
   wire FE_RN_517_0;
   wire FE_RN_516_0;
   wire FE_RN_515_0;
   wire FE_RN_514_0;
   wire FE_RN_513_0;
   wire FE_RN_512_0;
   wire FE_RN_511_0;
   wire FE_RN_510_0;
   wire FE_RN_509_0;
   wire FE_RN_477_0;
   wire FE_RN_476_0;
   wire FE_RN_475_0;
   wire FE_RN_474_0;
   wire FE_RN_473_0;
   wire FE_RN_472_0;
   wire FE_RN_471_0;
   wire FE_RN_470_0;
   wire FE_RN_469_0;
   wire FE_RN_468_0;
   wire FE_RN_467_0;
   wire FE_RN_466_0;
   wire FE_RN_465_0;
   wire FE_RN_464_0;
   wire FE_RN_463_0;
   wire FE_RN_462_0;
   wire FE_RN_461_0;
   wire FE_RN_460_0;
   wire FE_RN_459_0;
   wire FE_RN_458_0;
   wire FE_RN_457_0;
   wire FE_RN_456_0;
   wire FE_RN_455_0;
   wire FE_RN_454_0;
   wire FE_RN_453_0;
   wire FE_RN_434_0;
   wire FE_RN_433_0;
   wire FE_RN_432_0;
   wire FE_RN_431_0;
   wire FE_RN_430_0;
   wire FE_RN_429_0;
   wire FE_RN_428_0;
   wire FE_RN_427_0;
   wire FE_RN_426_0;
   wire FE_RN_425_0;
   wire FE_RN_424_0;
   wire FE_RN_423_0;
   wire FE_RN_422_0;
   wire FE_RN_421_0;
   wire FE_RN_420_0;
   wire FE_RN_419_0;
   wire FE_RN_418_0;
   wire FE_RN_417_0;
   wire FE_RN_416_0;
   wire FE_RN_415_0;
   wire FE_RN_414_0;
   wire FE_RN_413_0;
   wire FE_RN_383_0;
   wire FE_RN_382_0;
   wire FE_RN_381_0;
   wire FE_RN_380_0;
   wire FE_RN_375_0;
   wire FE_RN_374_0;
   wire FE_RN_373_0;
   wire FE_RN_372_0;
   wire FE_RN_371_0;
   wire FE_RN_370_0;
   wire FE_RN_369_0;
   wire FE_RN_368_0;
   wire FE_RN_367_0;
   wire FE_RN_366_0;
   wire FE_RN_365_0;
   wire FE_RN_364_0;
   wire FE_RN_363_0;
   wire FE_RN_362_0;
   wire FE_RN_361_0;
   wire FE_RN_360_0;
   wire FE_RN_359_0;
   wire FE_RN_358_0;
   wire FE_RN_357_0;
   wire FE_RN_356_0;
   wire FE_RN_355_0;
   wire FE_RN_354_0;
   wire FE_RN_353_0;
   wire FE_RN_352_0;
   wire FE_RN_351_0;
   wire FE_RN_350_0;
   wire FE_RN_349_0;
   wire FE_RN_348_0;
   wire FE_RN_347_0;
   wire FE_RN_346_0;
   wire FE_RN_345_0;
   wire FE_RN_344_0;
   wire FE_RN_343_0;
   wire FE_RN_342_0;
   wire FE_RN_341_0;
   wire FE_RN_340_0;
   wire FE_RN_339_0;
   wire FE_RN_338_0;
   wire FE_RN_337_0;
   wire FE_RN_336_0;
   wire FE_RN_335_0;
   wire FE_RN_334_0;
   wire FE_RN_333_0;
   wire FE_RN_332_0;
   wire FE_RN_331_0;
   wire FE_RN_330_0;
   wire FE_RN_329_0;
   wire FE_RN_328_0;
   wire FE_RN_327_0;
   wire FE_RN_326_0;
   wire FE_RN_325_0;
   wire FE_RN_324_0;
   wire FE_RN_322_0;
   wire FE_RN_321_0;
   wire FE_RN_320_0;
   wire FE_RN_319_0;
   wire FE_RN_318_0;
   wire FE_RN_317_0;
   wire FE_RN_316_0;
   wire FE_RN_315_0;
   wire FE_RN_314_0;
   wire FE_RN_313_0;
   wire FE_RN_312_0;
   wire FE_RN_311_0;
   wire FE_RN_310_0;
   wire FE_RN_309_0;
   wire FE_RN_308_0;
   wire FE_RN_307_0;
   wire FE_RN_306_0;
   wire FE_RN_305_0;
   wire FE_RN_304_0;
   wire FE_RN_303_0;
   wire FE_RN_302_0;
   wire FE_RN_301_0;
   wire FE_RN_300_0;
   wire FE_RN_299_0;
   wire FE_RN_298_0;
   wire FE_RN_276_0;
   wire FE_RN_275_0;
   wire FE_RN_274_0;
   wire FE_RN_273_0;
   wire FE_RN_272_0;
   wire FE_RN_270_0;
   wire FE_RN_269_0;
   wire FE_RN_268_0;
   wire FE_RN_266_0;
   wire FE_RN_265_0;
   wire FE_RN_264_0;
   wire FE_RN_263_0;
   wire FE_RN_262_0;
   wire FE_RN_261_0;
   wire FE_RN_260_0;
   wire FE_RN_259_0;
   wire FE_RN_258_0;
   wire FE_RN_257_0;
   wire FE_RN_256_0;
   wire FE_RN_254_0;
   wire FE_RN_253_0;
   wire FE_RN_252_0;
   wire FE_RN_251_0;
   wire FE_RN_250_0;
   wire FE_RN_249_0;
   wire FE_RN_248_0;
   wire FE_RN_247_0;
   wire FE_RN_246_0;
   wire FE_RN_245_0;
   wire FE_RN_244_0;
   wire FE_RN_242_0;
   wire FE_RN_241_0;
   wire FE_RN_240_0;
   wire FE_RN_239_0;
   wire FE_RN_238_0;
   wire FE_RN_237_0;
   wire FE_RN_236_0;
   wire FE_RN_235_0;
   wire FE_RN_234_0;
   wire FE_RN_233_0;
   wire FE_RN_232_0;
   wire FE_RN_231_0;
   wire FE_RN_230_0;
   wire FE_RN_229_0;
   wire FE_RN_228_0;
   wire FE_RN_227_0;
   wire FE_RN_226_0;
   wire FE_RN_225_0;
   wire FE_RN_224_0;
   wire FE_RN_223_0;
   wire FE_RN_222_0;
   wire FE_RN_192_0;
   wire FE_RN_191_0;
   wire FE_RN_190_0;
   wire FE_RN_189_0;
   wire FE_RN_187_0;
   wire FE_RN_182_0;
   wire FE_RN_181_0;
   wire FE_RN_180_0;
   wire FE_RN_179_0;
   wire FE_RN_178_0;
   wire FE_RN_177_0;
   wire FE_RN_176_0;
   wire FE_RN_175_0;
   wire FE_RN_174_0;
   wire FE_RN_173_0;
   wire FE_RN_172_0;
   wire FE_RN_171_0;
   wire FE_RN_170_0;
   wire FE_RN_169_0;
   wire FE_RN_168_0;
   wire FE_RN_167_0;
   wire FE_RN_166_0;
   wire FE_RN_165_0;
   wire FE_RN_164_0;
   wire FE_RN_163_0;
   wire FE_RN_162_0;
   wire FE_RN_161_0;
   wire FE_RN_160_0;
   wire FE_RN_159_0;
   wire FE_RN_158_0;
   wire FE_RN_157_0;
   wire FE_RN_156_0;
   wire FE_RN_155_0;
   wire FE_RN_154_0;
   wire FE_RN_153_0;
   wire FE_RN_152_0;
   wire FE_RN_151_0;
   wire FE_RN_150_0;
   wire FE_RN_149_0;
   wire FE_RN_148_0;
   wire FE_RN_147_0;
   wire FE_RN_146_0;
   wire FE_RN_145_0;
   wire FE_RN_144_0;
   wire FE_RN_143_0;
   wire FE_RN_142_0;
   wire FE_RN_141_0;
   wire FE_RN_140_0;
   wire FE_RN_139_0;
   wire FE_RN_138_0;
   wire FE_RN_137_0;
   wire FE_RN_136_0;
   wire FE_RN_135_0;
   wire FE_RN_134_0;
   wire FE_RN_133_0;
   wire FE_RN_132_0;
   wire FE_RN_131_0;
   wire FE_RN_130_0;
   wire FE_RN_129_0;
   wire FE_RN_128_0;
   wire FE_RN_127_0;
   wire FE_RN_126_0;
   wire FE_RN_125_0;
   wire FE_RN_124_0;
   wire FE_RN_123_0;
   wire FE_RN_122_0;
   wire FE_RN_121_0;
   wire FE_RN_120_0;
   wire FE_RN_119_0;
   wire FE_RN_118_0;
   wire FE_RN_117_0;
   wire FE_RN_116_0;
   wire FE_RN_115_0;
   wire FE_RN_114_0;
   wire FE_RN_113_0;
   wire FE_RN_112_0;
   wire FE_RN_111_0;
   wire FE_RN_110_0;
   wire FE_RN_109_0;
   wire FE_RN_108_0;
   wire FE_RN_107_0;
   wire FE_RN_106_0;
   wire FE_RN_105_0;
   wire FE_RN_104_0;
   wire FE_RN_103_0;
   wire FE_RN_102_0;
   wire FE_RN_101_0;
   wire FE_RN_99_0;
   wire FE_RN_84_0;
   wire FE_RN_83_0;
   wire FE_RN_82_0;
   wire FE_RN_81_0;
   wire FE_RN_80_0;
   wire FE_RN_79_0;
   wire FE_RN_78_0;
   wire FE_RN_77_0;
   wire FE_RN_76_0;
   wire FE_RN_75_0;
   wire FE_RN_74_0;
   wire FE_RN_73_0;
   wire FE_RN_72_0;
   wire FE_RN_71_0;
   wire FE_RN_70_0;
   wire FE_RN_69_0;
   wire FE_RN_68_0;
   wire FE_RN_67_0;
   wire FE_RN_66_0;
   wire FE_RN_65_0;
   wire FE_RN_64_0;
   wire FE_RN_63_0;
   wire FE_RN_62_0;
   wire FE_RN_61_0;
   wire FE_RN_60_0;
   wire FE_RN_59_0;
   wire FE_RN_58_0;
   wire FE_RN_57_0;
   wire FE_RN_56_0;
   wire FE_RN_55_0;
   wire FE_RN_54_0;
   wire FE_RN_53_0;
   wire FE_RN_52_0;
   wire FE_RN_51_0;
   wire FE_RN_50_0;
   wire FE_RN_49_0;
   wire FE_RN_48_0;
   wire FE_RN_47_0;
   wire FE_RN_46_0;
   wire FE_RN_45_0;
   wire FE_RN_44_0;
   wire FE_RN_43_0;
   wire FE_RN_42_0;
   wire FE_RN_41_0;
   wire FE_RN_40_0;
   wire FE_RN_39_0;
   wire FE_RN_38_0;
   wire FE_RN_37_0;
   wire FE_RN_36_0;
   wire FE_RN_35_0;
   wire FE_RN_34_0;
   wire FE_RN_31_0;
   wire FE_RN_30_0;
   wire FE_RN_29_0;
   wire FE_RN_28_0;
   wire FE_RN_27_0;
   wire FE_RN_26_0;
   wire FE_RN_25_0;
   wire FE_RN_24_0;
   wire FE_RN_23_0;
   wire FE_RN_22_0;
   wire FE_RN_20_0;
   wire FE_RN_19_0;
   wire FE_RN_18_0;
   wire FE_RN_16_0;
   wire FE_RN_15_0;
   wire FE_RN_14_0;
   wire FE_RN_13_0;
   wire FE_RN_12_0;
   wire FE_RN_11_0;
   wire FE_RN_5_0;
   wire FE_RN_4_0;
   wire FE_RN_3_0;
   wire FE_RN_1_0;
   wire FE_RN_0_0;
   wire \u_div/SumTmp[1][0] ;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][3] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[5][3] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;

   CLKNAND2X2M FE_RC_651_0 (.Y(FE_RN_543_0), 
	.B(FE_RN_517_0), 
	.A(FE_RN_519_0));
   NAND3BX4M FE_RC_650_0 (.Y(FE_RN_509_0), 
	.C(FE_RN_515_0), 
	.B(FE_RN_510_0), 
	.AN(FE_RN_543_0));
   INVX2M FE_RC_649_0 (.Y(FE_RN_542_0), 
	.A(FE_RN_515_0));
   INVX2M FE_RC_648_0 (.Y(FE_RN_541_0), 
	.A(FE_RN_540_0));
   NAND2X4M FE_RC_647_0 (.Y(FE_RN_540_0), 
	.B(FE_RN_520_0), 
	.A(FE_RN_521_0));
   INVX2M FE_RC_646_0 (.Y(FE_RN_539_0), 
	.A(FE_RN_522_0));
   AOI2B1X4M FE_RC_645_0 (.Y(FE_RN_538_0), 
	.B0(FE_RN_539_0), 
	.A1N(FE_RN_519_0), 
	.A0(FE_RN_540_0));
   OAI2B1X4M FE_RC_644_0 (.Y(FE_RN_537_0), 
	.B0(FE_RN_538_0), 
	.A1N(FE_RN_540_0), 
	.A0(FE_RN_517_0));
   AOI2B1X4M FE_RC_643_0 (.Y(FE_RN_536_0), 
	.B0(FE_RN_537_0), 
	.A1N(FE_RN_541_0), 
	.A0(FE_RN_542_0));
   OAI2B1X4M FE_RC_642_0 (.Y(FE_RN_535_0), 
	.B0(FE_RN_536_0), 
	.A1N(FE_RN_540_0), 
	.A0(FE_RN_510_0));
   AND2X8M FE_RC_641_0 (.Y(quotient[1]), 
	.B(n12), 
	.A(FE_RN_535_0));
   INVX2M FE_RC_640_0 (.Y(FE_RN_534_0), 
	.A(FE_RN_519_0));
   NOR2X4M FE_RC_639_0 (.Y(FE_RN_533_0), 
	.B(FE_RN_534_0), 
	.A(FE_RN_523_0));
   INVX2M FE_RC_638_0 (.Y(FE_RN_532_0), 
	.A(FE_RN_511_0));
   OAI21X4M FE_RC_637_0 (.Y(FE_RN_531_0), 
	.B0(FE_RN_530_0), 
	.A1(FE_RN_532_0), 
	.A0(FE_RN_533_0));
   XOR2X2M FE_RC_636_0 (.Y(FE_RN_530_0), 
	.B(n173), 
	.A(\u_div/PartRem[2][6] ));
   INVX2M FE_RC_635_0 (.Y(FE_RN_529_0), 
	.A(FE_RN_530_0));
   NAND2X4M FE_RC_634_0 (.Y(FE_RN_528_0), 
	.B(FE_RN_529_0), 
	.A(FE_RN_509_0));
   NAND2X3M FE_RC_633_0 (.Y(\u_div/SumTmp[1][6] ), 
	.B(FE_RN_531_0), 
	.A(FE_RN_528_0));
   XNOR2X2M FE_RC_632_0 (.Y(FE_RN_527_0), 
	.B(n14), 
	.A(\u_div/PartRem[2][5] ));
   INVX2M FE_RC_631_0 (.Y(FE_RN_526_0), 
	.A(FE_RN_511_0));
   NOR2BX2M FE_RC_630_0 (.Y(FE_RN_525_0), 
	.B(FE_RN_526_0), 
	.AN(FE_RN_519_0));
   INVX2M FE_RC_629_0 (.Y(FE_RN_524_0), 
	.A(FE_RN_462_0));
   NAND3BX4M FE_RC_628_0 (.Y(FE_RN_523_0), 
	.C(FE_RN_459_0), 
	.B(FE_RN_453_0), 
	.AN(FE_RN_524_0));
   MXI2X2M FE_RC_627_0 (.Y(\u_div/SumTmp[1][5] ), 
	.S0(FE_RN_523_0), 
	.B(FE_RN_525_0), 
	.A(FE_RN_527_0));
   CLKNAND2X2M FE_RC_626_0 (.Y(FE_RN_522_0), 
	.B(n173), 
	.A(\u_div/PartRem[2][6] ));
   INVX2M FE_RC_625_0 (.Y(FE_RN_521_0), 
	.A(n173));
   INVX2M FE_RC_624_0 (.Y(FE_RN_520_0), 
	.A(\u_div/PartRem[2][6] ));
   CLKNAND2X4M FE_RC_623_0 (.Y(FE_RN_519_0), 
	.B(n14), 
	.A(\u_div/PartRem[2][5] ));
   INVX2M FE_RC_622_0 (.Y(FE_RN_518_0), 
	.A(FE_RN_462_0));
   CLKNAND2X4M FE_RC_621_0 (.Y(FE_RN_517_0), 
	.B(FE_RN_518_0), 
	.A(FE_RN_511_0));
   INVX2M FE_RC_620_0 (.Y(FE_RN_516_0), 
	.A(FE_RN_459_0));
   CLKNAND2X4M FE_RC_619_0 (.Y(FE_RN_515_0), 
	.B(FE_RN_516_0), 
	.A(FE_RN_511_0));
   INVX2M FE_RC_618_0 (.Y(FE_RN_514_0), 
	.A(FE_RN_453_0));
   INVX2M FE_RC_617_0 (.Y(FE_RN_513_0), 
	.A(n14));
   INVX2M FE_RC_616_0 (.Y(FE_RN_512_0), 
	.A(\u_div/PartRem[2][5] ));
   NAND2X5M FE_RC_615_0 (.Y(FE_RN_511_0), 
	.B(FE_RN_513_0), 
	.A(FE_RN_512_0));
   NAND2X2M FE_RC_614_0 (.Y(FE_RN_510_0), 
	.B(FE_RN_514_0), 
	.A(FE_RN_511_0));
   XOR2X2M FE_RC_575_0 (.Y(FE_RN_477_0), 
	.B(n15), 
	.A(\u_div/PartRem[2][4] ));
   INVX2M FE_RC_574_0 (.Y(FE_RN_476_0), 
	.A(\u_div/CryTmp[1][3] ));
   NAND2X3M FE_RC_573_0 (.Y(FE_RN_475_0), 
	.B(FE_RN_476_0), 
	.A(FE_RN_461_0));
   NAND2X3M FE_RC_572_0 (.Y(FE_RN_474_0), 
	.B(FE_RN_454_0), 
	.A(FE_RN_475_0));
   NAND2X3M FE_RC_571_0 (.Y(FE_RN_473_0), 
	.B(FE_RN_477_0), 
	.A(FE_RN_474_0));
   INVX2M FE_RC_570_0 (.Y(FE_RN_472_0), 
	.A(FE_RN_461_0));
   NAND2X4M FE_RC_569_0 (.Y(FE_RN_471_0), 
	.B(FE_RN_472_0), 
	.A(FE_RN_469_0));
   CLKNAND2X2M FE_RC_568_0 (.Y(FE_RN_470_0), 
	.B(n15), 
	.A(\u_div/PartRem[2][4] ));
   CLKNAND2X4M FE_RC_567_0 (.Y(FE_RN_469_0), 
	.B(FE_RN_470_0), 
	.A(FE_RN_456_0));
   NAND3X4M FE_RC_566_0 (.Y(FE_RN_468_0), 
	.C(\u_div/CryTmp[1][3] ), 
	.B(FE_RN_454_0), 
	.A(FE_RN_469_0));
   NAND3X4M FE_RC_565_0 (.Y(\u_div/SumTmp[1][4] ), 
	.C(FE_RN_473_0), 
	.B(FE_RN_471_0), 
	.A(FE_RN_468_0));
   INVX2M FE_RC_564_0 (.Y(FE_RN_467_0), 
	.A(\u_div/CryTmp[1][3] ));
   XOR2X2M FE_RC_563_0 (.Y(FE_RN_466_0), 
	.B(n16), 
	.A(\u_div/PartRem[2][3] ));
   NAND2X2M FE_RC_562_0 (.Y(FE_RN_465_0), 
	.B(FE_RN_467_0), 
	.A(FE_RN_466_0));
   CLKNAND2X4M FE_RC_561_0 (.Y(FE_RN_464_0), 
	.B(FE_RN_461_0), 
	.A(FE_RN_454_0));
   NAND2X4M FE_RC_560_0 (.Y(FE_RN_463_0), 
	.B(\u_div/CryTmp[1][3] ), 
	.A(FE_RN_464_0));
   CLKNAND2X4M FE_RC_559_0 (.Y(\u_div/SumTmp[1][3] ), 
	.B(FE_RN_465_0), 
	.A(FE_RN_463_0));
   CLKNAND2X2M FE_RC_558_0 (.Y(FE_RN_462_0), 
	.B(n15), 
	.A(\u_div/PartRem[2][4] ));
   CLKNAND2X4M FE_RC_557_0 (.Y(FE_RN_461_0), 
	.B(n16), 
	.A(\u_div/PartRem[2][3] ));
   INVX2M FE_RC_556_0 (.Y(FE_RN_460_0), 
	.A(FE_RN_461_0));
   NAND2X4M FE_RC_555_0 (.Y(FE_RN_459_0), 
	.B(FE_RN_460_0), 
	.A(FE_RN_456_0));
   INVX2M FE_RC_554_0 (.Y(FE_RN_458_0), 
	.A(n15));
   INVX2M FE_RC_553_0 (.Y(FE_RN_457_0), 
	.A(\u_div/PartRem[2][4] ));
   NAND2X4M FE_RC_552_0 (.Y(FE_RN_456_0), 
	.B(FE_RN_458_0), 
	.A(FE_RN_457_0));
   INVX2M FE_RC_551_0 (.Y(FE_RN_455_0), 
	.A(n16));
   NAND2BX4M FE_RC_550_0 (.Y(FE_RN_454_0), 
	.B(FE_RN_455_0), 
	.AN(\u_div/PartRem[2][3] ));
   NAND3X4M FE_RC_549_0 (.Y(FE_RN_453_0), 
	.C(\u_div/CryTmp[1][3] ), 
	.B(FE_RN_456_0), 
	.A(FE_RN_454_0));
   INVX2M FE_RC_525_0 (.Y(FE_RN_434_0), 
	.A(\u_div/PartRem[3][1] ));
   INVX2M FE_RC_524_0 (.Y(FE_RN_433_0), 
	.A(\u_div/SumTmp[2][1] ));
   MXI2X6M FE_RC_523_0 (.Y(\u_div/PartRem[2][2] ), 
	.S0(quotient[2]), 
	.B(FE_RN_433_0), 
	.A(FE_RN_434_0));
   OAI2B1X4M FE_RC_522_0 (.Y(FE_RN_432_0), 
	.B0(FE_RN_416_0), 
	.A1N(FE_RN_418_0), 
	.A0(\u_div/PartRem[2][1] ));
   NAND2X4M FE_RC_521_0 (.Y(FE_RN_431_0), 
	.B(n17), 
	.A(FE_RN_421_0));
   CLKNAND2X4M FE_RC_520_0 (.Y(FE_RN_430_0), 
	.B(FE_RN_419_0), 
	.A(FE_RN_431_0));
   CLKNAND2X4M FE_RC_519_0 (.Y(FE_RN_429_0), 
	.B(FE_RN_430_0), 
	.A(FE_RN_414_0));
   OAI2B1X4M FE_RC_518_0 (.Y(\u_div/SumTmp[1][2] ), 
	.B0(FE_RN_429_0), 
	.A1N(FE_RN_432_0), 
	.A0(FE_RN_430_0));
   OAI2BB2X4M FE_RC_517_0 (.Y(FE_RN_428_0), 
	.B1(\u_div/CryTmp[1][1] ), 
	.B0(n18), 
	.A1N(n18), 
	.A0N(\u_div/CryTmp[1][1] ));
   NAND2X4M FE_RC_516_0 (.Y(FE_RN_427_0), 
	.B(FE_RN_418_0), 
	.A(FE_RN_416_0));
   NAND2X4M FE_RC_515_0 (.Y(FE_RN_426_0), 
	.B(\u_div/PartRem[2][1] ), 
	.A(FE_RN_427_0));
   OAI21X4M FE_RC_514_0 (.Y(\u_div/SumTmp[1][1] ), 
	.B0(FE_RN_426_0), 
	.A1(\u_div/PartRem[2][1] ), 
	.A0(FE_RN_428_0));
   NAND2X4M FE_RC_513_0 (.Y(FE_RN_425_0), 
	.B(n17), 
	.A(FE_RN_421_0));
   INVX2M FE_RC_512_0 (.Y(FE_RN_424_0), 
	.A(n17));
   INVX2M FE_RC_511_0 (.Y(FE_RN_423_0), 
	.A(\u_div/PartRem[3][1] ));
   INVX2M FE_RC_510_0 (.Y(FE_RN_422_0), 
	.A(\u_div/SumTmp[2][1] ));
   MXI2X6M FE_RC_509_0 (.Y(FE_RN_421_0), 
	.S0(quotient[2]), 
	.B(FE_RN_422_0), 
	.A(FE_RN_423_0));
   INVX2M FE_RC_508_0 (.Y(FE_RN_420_0), 
	.A(FE_RN_421_0));
   NAND2X3M FE_RC_507_0 (.Y(FE_RN_419_0), 
	.B(FE_RN_424_0), 
	.A(FE_RN_420_0));
   NAND2X4M FE_RC_506_0 (.Y(FE_RN_418_0), 
	.B(\u_div/CryTmp[1][1] ), 
	.A(n18));
   INVX2M FE_RC_505_0 (.Y(FE_RN_417_0), 
	.A(n18));
   NAND2BX8M FE_RC_504_0 (.Y(FE_RN_416_0), 
	.B(FE_RN_417_0), 
	.AN(\u_div/CryTmp[1][1] ));
   NAND2X4M FE_RC_503_0 (.Y(FE_RN_415_0), 
	.B(\u_div/PartRem[2][1] ), 
	.A(FE_RN_416_0));
   CLKNAND2X4M FE_RC_502_0 (.Y(FE_RN_414_0), 
	.B(FE_RN_418_0), 
	.A(FE_RN_415_0));
   CLKNAND2X4M FE_RC_501_0 (.Y(FE_RN_413_0), 
	.B(FE_RN_419_0), 
	.A(FE_RN_414_0));
   NAND2X3M FE_RC_500_0 (.Y(\u_div/CryTmp[1][3] ), 
	.B(FE_RN_425_0), 
	.A(FE_RN_413_0));
   AND2X8M FE_RC_467_0 (.Y(quotient[2]), 
	.B(n22), 
	.A(\u_div/CryTmp[2][6] ));
   INVX2M FE_RC_466_0 (.Y(FE_RN_383_0), 
	.A(n22));
   NAND3BX4M FE_RC_465_0 (.Y(FE_RN_382_0), 
	.C(\u_div/SumTmp[2][0] ), 
	.B(\u_div/CryTmp[2][6] ), 
	.AN(FE_RN_383_0));
   INVX2M FE_RC_464_0 (.Y(FE_RN_381_0), 
	.A(n22));
   CLKNAND2X4M FE_RC_463_0 (.Y(FE_RN_380_0), 
	.B(FE_RN_381_0), 
	.A(a[2]));
   OAI2B11X4M FE_RC_462_0 (.Y(\u_div/PartRem[2][1] ), 
	.C0(FE_RN_380_0), 
	.B0(FE_RN_382_0), 
	.A1N(a[2]), 
	.A0(\u_div/CryTmp[2][6] ));
   INVX2M FE_RC_455_0 (.Y(FE_RN_375_0), 
	.A(n14));
   INVX2M FE_RC_454_0 (.Y(FE_RN_374_0), 
	.A(\u_div/PartRem[3][5] ));
   INVX2M FE_RC_453_0 (.Y(FE_RN_373_0), 
	.A(FE_RN_359_0));
   OAI2BB1X2M FE_RC_452_0 (.Y(FE_RN_372_0), 
	.B0(FE_RN_373_0), 
	.A1N(FE_RN_374_0), 
	.A0N(FE_RN_375_0));
   INVX2M FE_RC_451_0 (.Y(FE_RN_371_0), 
	.A(FE_RN_336_0));
   NAND4BBX4M FE_RC_450_0 (.Y(FE_RN_370_0), 
	.D(FE_RN_362_0), 
	.C(FE_RN_338_0), 
	.BN(FE_RN_371_0), 
	.AN(FE_RN_372_0));
   INVX2M FE_RC_449_0 (.Y(FE_RN_369_0), 
	.A(FE_RN_359_0));
   NAND2X3M FE_RC_448_0 (.Y(FE_RN_368_0), 
	.B(FE_RN_364_0), 
	.A(FE_RN_369_0));
   CLKNAND2X4M FE_RC_447_0 (.Y(FE_RN_367_0), 
	.B(FE_RN_368_0), 
	.A(FE_RN_361_0));
   OAI2B11X2M FE_RC_446_0 (.Y(\u_div/SumTmp[2][5] ), 
	.C0(FE_RN_367_0), 
	.B0(FE_RN_370_0), 
	.A1N(FE_RN_368_0), 
	.A0(FE_RN_338_0));
   INVX2M FE_RC_445_0 (.Y(FE_RN_366_0), 
	.A(n14));
   INVX2M FE_RC_444_0 (.Y(FE_RN_365_0), 
	.A(\u_div/PartRem[3][5] ));
   NAND2X2M FE_RC_443_0 (.Y(FE_RN_364_0), 
	.B(FE_RN_366_0), 
	.A(FE_RN_365_0));
   INVX2M FE_RC_442_0 (.Y(FE_RN_363_0), 
	.A(FE_RN_327_0));
   NAND2X4M FE_RC_441_0 (.Y(FE_RN_362_0), 
	.B(FE_RN_339_0), 
	.A(FE_RN_363_0));
   NAND2X4M FE_RC_440_0 (.Y(FE_RN_361_0), 
	.B(FE_RN_336_0), 
	.A(FE_RN_362_0));
   CLKNAND2X4M FE_RC_439_0 (.Y(FE_RN_360_0), 
	.B(FE_RN_364_0), 
	.A(FE_RN_361_0));
   AND2X2M FE_RC_438_0 (.Y(FE_RN_359_0), 
	.B(n14), 
	.A(\u_div/PartRem[3][5] ));
   INVX2M FE_RC_437_0 (.Y(FE_RN_358_0), 
	.A(FE_RN_359_0));
   OAI2B11X4M FE_RC_436_0 (.Y(\u_div/CryTmp[2][6] ), 
	.C0(FE_RN_358_0), 
	.B0(FE_RN_360_0), 
	.A1N(FE_RN_364_0), 
	.A0(FE_RN_338_0));
   INVX2M FE_RC_435_0 (.Y(FE_RN_357_0), 
	.A(FE_RN_327_0));
   CLKNAND2X4M FE_RC_434_0 (.Y(FE_RN_356_0), 
	.B(FE_RN_357_0), 
	.A(FE_RN_354_0));
   INVX2M FE_RC_433_0 (.Y(FE_RN_355_0), 
	.A(FE_RN_337_0));
   NAND2X3M FE_RC_432_0 (.Y(FE_RN_354_0), 
	.B(FE_RN_339_0), 
	.A(FE_RN_355_0));
   NAND3X4M FE_RC_431_0 (.Y(FE_RN_353_0), 
	.C(FE_RN_325_0), 
	.B(FE_RN_324_0), 
	.A(FE_RN_354_0));
   INVX2M FE_RC_430_0 (.Y(FE_RN_352_0), 
	.A(FE_RN_324_0));
   INVX2M FE_RC_429_0 (.Y(FE_RN_351_0), 
	.A(FE_RN_344_0));
   NAND3X3M FE_RC_428_0 (.Y(FE_RN_350_0), 
	.C(FE_RN_327_0), 
	.B(FE_RN_352_0), 
	.A(FE_RN_351_0));
   INVX2M FE_RC_427_0 (.Y(FE_RN_349_0), 
	.A(FE_RN_325_0));
   INVX2M FE_RC_426_0 (.Y(FE_RN_348_0), 
	.A(n15));
   INVX2M FE_RC_425_0 (.Y(FE_RN_347_0), 
	.A(\u_div/PartRem[3][4] ));
   NAND2X2M FE_RC_424_0 (.Y(FE_RN_346_0), 
	.B(FE_RN_348_0), 
	.A(FE_RN_347_0));
   INVX2M FE_RC_423_0 (.Y(FE_RN_345_0), 
	.A(FE_RN_337_0));
   NAND2X3M FE_RC_422_0 (.Y(FE_RN_344_0), 
	.B(FE_RN_346_0), 
	.A(FE_RN_345_0));
   INVX2M FE_RC_421_0 (.Y(FE_RN_343_0), 
	.A(FE_RN_344_0));
   NAND3X3M FE_RC_420_0 (.Y(FE_RN_342_0), 
	.C(FE_RN_327_0), 
	.B(FE_RN_349_0), 
	.A(FE_RN_343_0));
   NAND4X2M FE_RC_419_0 (.Y(\u_div/SumTmp[2][4] ), 
	.D(FE_RN_356_0), 
	.C(FE_RN_353_0), 
	.B(FE_RN_350_0), 
	.A(FE_RN_342_0));
   INVX2M FE_RC_418_0 (.Y(FE_RN_341_0), 
	.A(n15));
   INVX2M FE_RC_417_0 (.Y(FE_RN_340_0), 
	.A(\u_div/PartRem[3][4] ));
   NAND2X4M FE_RC_416_0 (.Y(FE_RN_339_0), 
	.B(FE_RN_341_0), 
	.A(FE_RN_340_0));
   NAND3X4M FE_RC_415_0 (.Y(FE_RN_338_0), 
	.C(FE_RN_325_0), 
	.B(FE_RN_324_0), 
	.A(FE_RN_339_0));
   CLKAND2X6M FE_RC_414_0 (.Y(FE_RN_337_0), 
	.B(n15), 
	.A(\u_div/PartRem[3][4] ));
   INVX2M FE_RC_413_0 (.Y(FE_RN_336_0), 
	.A(FE_RN_337_0));
   INVX2M FE_RC_411_0 (.Y(FE_RN_335_0), 
	.A(n16));
   INVX2M FE_RC_410_0 (.Y(FE_RN_334_0), 
	.A(\u_div/PartRem[3][3] ));
   INVX2M FE_RC_409_0 (.Y(FE_RN_333_0), 
	.A(FE_RN_328_0));
   OAI2BB1X2M FE_RC_408_0 (.Y(FE_RN_332_0), 
	.B0(FE_RN_333_0), 
	.A1N(FE_RN_334_0), 
	.A0N(FE_RN_335_0));
   INVX2M FE_RC_407_0 (.Y(FE_RN_331_0), 
	.A(FE_RN_325_0));
   NOR2X2M FE_RC_406_0 (.Y(FE_RN_330_0), 
	.B(FE_RN_331_0), 
	.A(FE_RN_328_0));
   MXI2X2M FE_RC_405_0 (.Y(\u_div/SumTmp[2][3] ), 
	.S0(FE_RN_324_0), 
	.B(FE_RN_330_0), 
	.A(FE_RN_332_0));
   INVX2M FE_RC_404_0 (.Y(FE_RN_329_0), 
	.A(n16));
   NOR2BX4M FE_RC_403_0 (.Y(FE_RN_328_0), 
	.B(FE_RN_329_0), 
	.AN(\u_div/PartRem[3][3] ));
   INVX2M FE_RC_402_0 (.Y(FE_RN_327_0), 
	.A(FE_RN_328_0));
   INVX2M FE_RC_401_0 (.Y(FE_RN_326_0), 
	.A(n16));
   NAND2BX4M FE_RC_400_0 (.Y(FE_RN_325_0), 
	.B(FE_RN_326_0), 
	.AN(\u_div/PartRem[3][3] ));
   NAND2X6M FE_RC_399_0 (.Y(FE_RN_324_0), 
	.B(FE_RN_307_0), 
	.A(FE_RN_298_0));
   CLKNAND2X4M FE_RC_396_0 (.Y(FE_RN_272_0), 
	.B(FE_RN_273_0), 
	.A(FE_RN_256_0));
   MXI2X4M FE_RC_395_0 (.Y(\u_div/PartRem[3][1] ), 
	.S0(FE_RN_304_0), 
	.B(FE_RN_275_0), 
	.A(FE_RN_276_0));
   INVX2M FE_RC_394_0 (.Y(FE_RN_322_0), 
	.A(FE_RN_299_0));
   INVX2M FE_RC_393_0 (.Y(FE_RN_321_0), 
	.A(\u_div/CryTmp[2][1] ));
   INVX2M FE_RC_392_0 (.Y(FE_RN_320_0), 
	.A(FE_RN_301_0));
   AOI21X2M FE_RC_391_0 (.Y(FE_RN_319_0), 
	.B0(FE_RN_320_0), 
	.A1(FE_RN_321_0), 
	.A0(FE_RN_306_0));
   XOR2X4M FE_RC_390_0 (.Y(FE_RN_318_0), 
	.B(n17), 
	.A(\u_div/PartRem[3][2] ));
   MXI2X2M FE_RC_389_0 (.Y(\u_div/SumTmp[2][2] ), 
	.S0(FE_RN_318_0), 
	.B(FE_RN_319_0), 
	.A(FE_RN_322_0));
   CLKNAND2X8M FE_RC_388_0 (.Y(FE_RN_317_0), 
	.B(FE_RN_306_0), 
	.A(FE_RN_301_0));
   NAND2X3M FE_RC_387_0 (.Y(FE_RN_316_0), 
	.B(\u_div/CryTmp[2][1] ), 
	.A(FE_RN_317_0));
   INVX2M FE_RC_386_0 (.Y(FE_RN_315_0), 
	.A(\u_div/CryTmp[2][1] ));
   XNOR2X4M FE_RC_385_0 (.Y(FE_RN_314_0), 
	.B(n18), 
	.A(FE_RN_303_0));
   INVX2M FE_RC_384_0 (.Y(FE_RN_313_0), 
	.A(FE_RN_314_0));
   NAND2X3M FE_RC_383_0 (.Y(FE_RN_312_0), 
	.B(FE_RN_315_0), 
	.A(FE_RN_313_0));
   NAND2X2M FE_RC_382_0 (.Y(\u_div/SumTmp[2][1] ), 
	.B(FE_RN_316_0), 
	.A(FE_RN_312_0));
   INVX2M FE_RC_381_0 (.Y(FE_RN_311_0), 
	.A(n17));
   AND2X4M FE_RC_380_0 (.Y(FE_RN_310_0), 
	.B(FE_RN_311_0), 
	.A(FE_RN_306_0));
   CLKNAND2X8M FE_RC_379_0 (.Y(FE_RN_309_0), 
	.B(\u_div/CryTmp[2][1] ), 
	.A(FE_RN_301_0));
   NAND2X4M FE_RC_378_0 (.Y(FE_RN_308_0), 
	.B(FE_RN_310_0), 
	.A(FE_RN_309_0));
   NAND2X4M FE_RC_377_0 (.Y(FE_RN_307_0), 
	.B(\u_div/PartRem[3][2] ), 
	.A(FE_RN_308_0));
   NAND2X6M FE_RC_376_0 (.Y(FE_RN_306_0), 
	.B(n18), 
	.A(FE_RN_303_0));
   CLKNAND2X4M FE_RC_375_0 (.Y(FE_RN_305_0), 
	.B(FE_RN_256_0), 
	.A(FE_RN_273_0));
   NAND2X5M FE_RC_374_0 (.Y(FE_RN_304_0), 
	.B(FE_RN_269_0), 
	.A(FE_RN_305_0));
   MXI2X6M FE_RC_373_0 (.Y(FE_RN_303_0), 
	.S0(FE_RN_304_0), 
	.B(FE_RN_275_0), 
	.A(FE_RN_276_0));
   INVX2M FE_RC_372_0 (.Y(FE_RN_302_0), 
	.A(n18));
   NAND2BX8M FE_RC_371_0 (.Y(FE_RN_301_0), 
	.B(FE_RN_302_0), 
	.AN(FE_RN_303_0));
   CLKNAND2X8M FE_RC_370_0 (.Y(FE_RN_300_0), 
	.B(\u_div/CryTmp[2][1] ), 
	.A(FE_RN_301_0));
   NAND2X4M FE_RC_369_0 (.Y(FE_RN_299_0), 
	.B(FE_RN_306_0), 
	.A(FE_RN_300_0));
   NAND2X4M FE_RC_368_0 (.Y(FE_RN_298_0), 
	.B(n17), 
	.A(FE_RN_299_0));
   NAND2X6M FE_RC_340_0 (.Y(quotient[3]), 
	.B(FE_RN_272_0), 
	.A(FE_RN_269_0));
   INVX2M FE_RC_339_0 (.Y(FE_RN_276_0), 
	.A(a[3]));
   INVX2M FE_RC_338_0 (.Y(FE_RN_275_0), 
	.A(\u_div/SumTmp[3][0] ));
   INVX2M FE_RC_337_0 (.Y(FE_RN_274_0), 
	.A(FE_RN_268_0));
   NOR2BX4M FE_RC_336_0 (.Y(FE_RN_273_0), 
	.B(FE_RN_274_0), 
	.AN(FE_RN_258_0));
   AND2X2M FE_RC_332_0 (.Y(FE_RN_270_0), 
	.B(n14), 
	.A(n22));
   NAND2BX4M FE_RC_331_0 (.Y(FE_RN_269_0), 
	.B(FE_RN_270_0), 
	.AN(FE_RN_259_0));
   AND2X2M FE_RC_330_0 (.Y(FE_RN_268_0), 
	.B(n14), 
	.A(n22));
   INVX2M FE_RC_327_0 (.Y(FE_RN_266_0), 
	.A(n15));
   INVX2M FE_RC_326_0 (.Y(FE_RN_265_0), 
	.A(\u_div/PartRem[4][4] ));
   INVX2M FE_RC_325_0 (.Y(FE_RN_264_0), 
	.A(FE_RN_260_0));
   OAI2BB1X2M FE_RC_324_0 (.Y(FE_RN_263_0), 
	.B0(FE_RN_264_0), 
	.A1N(FE_RN_265_0), 
	.A0N(FE_RN_266_0));
   INVX2M FE_RC_323_0 (.Y(FE_RN_262_0), 
	.A(FE_RN_258_0));
   NOR2X4M FE_RC_322_0 (.Y(FE_RN_261_0), 
	.B(FE_RN_262_0), 
	.A(FE_RN_260_0));
   MXI2X2M FE_RC_321_0 (.Y(\u_div/SumTmp[3][4] ), 
	.S0(FE_RN_256_0), 
	.B(FE_RN_261_0), 
	.A(FE_RN_263_0));
   AND2X2M FE_RC_320_0 (.Y(FE_RN_260_0), 
	.B(n15), 
	.A(\u_div/PartRem[4][4] ));
   INVX2M FE_RC_319_0 (.Y(FE_RN_259_0), 
	.A(FE_RN_260_0));
   OR2X2M FE_RC_318_0 (.Y(FE_RN_258_0), 
	.B(n15), 
	.A(\u_div/PartRem[4][4] ));
   NAND2X4M FE_RC_317_0 (.Y(FE_RN_257_0), 
	.B(FE_RN_245_0), 
	.A(FE_RN_244_0));
   NAND2X6M FE_RC_316_0 (.Y(FE_RN_256_0), 
	.B(FE_RN_247_0), 
	.A(FE_RN_257_0));
   INVX2M FE_RC_313_0 (.Y(FE_RN_254_0), 
	.A(n16));
   INVX2M FE_RC_312_0 (.Y(FE_RN_253_0), 
	.A(\u_div/PartRem[4][3] ));
   INVX2M FE_RC_311_0 (.Y(FE_RN_252_0), 
	.A(FE_RN_248_0));
   OAI2BB1X2M FE_RC_310_0 (.Y(FE_RN_251_0), 
	.B0(FE_RN_252_0), 
	.A1N(FE_RN_253_0), 
	.A0N(FE_RN_254_0));
   INVX2M FE_RC_309_0 (.Y(FE_RN_250_0), 
	.A(FE_RN_245_0));
   NOR2X4M FE_RC_308_0 (.Y(FE_RN_249_0), 
	.B(FE_RN_250_0), 
	.A(FE_RN_248_0));
   MXI2X1M FE_RC_307_0 (.Y(\u_div/SumTmp[3][3] ), 
	.S0(FE_RN_244_0), 
	.B(FE_RN_249_0), 
	.A(FE_RN_251_0));
   CLKAND2X4M FE_RC_306_0 (.Y(FE_RN_248_0), 
	.B(n16), 
	.A(\u_div/PartRem[4][3] ));
   INVX2M FE_RC_305_0 (.Y(FE_RN_247_0), 
	.A(FE_RN_248_0));
   INVX2M FE_RC_304_0 (.Y(FE_RN_246_0), 
	.A(\u_div/PartRem[4][3] ));
   NAND2BX2M FE_RC_303_0 (.Y(FE_RN_245_0), 
	.B(FE_RN_246_0), 
	.AN(n16));
   NAND2X6M FE_RC_302_0 (.Y(FE_RN_244_0), 
	.B(FE_RN_231_0), 
	.A(FE_RN_222_0));
   NAND2X4M FE_RC_299_0 (.Y(FE_RN_187_0), 
	.B(FE_RN_229_0), 
	.A(n21));
   MXI2X4M FE_RC_298_0 (.Y(\u_div/PartRem[4][1] ), 
	.S0(FE_RN_228_0), 
	.B(FE_RN_191_0), 
	.A(FE_RN_192_0));
   INVX2M FE_RC_297_0 (.Y(FE_RN_242_0), 
	.A(FE_RN_223_0));
   INVX2M FE_RC_296_0 (.Y(FE_RN_241_0), 
	.A(\u_div/CryTmp[3][1] ));
   INVX2M FE_RC_295_0 (.Y(FE_RN_240_0), 
	.A(FE_RN_225_0));
   AOI21X4M FE_RC_294_0 (.Y(FE_RN_239_0), 
	.B0(FE_RN_240_0), 
	.A1(FE_RN_241_0), 
	.A0(FE_RN_230_0));
   XOR2X4M FE_RC_293_0 (.Y(FE_RN_238_0), 
	.B(n17), 
	.A(\u_div/PartRem[4][2] ));
   MXI2X2M FE_RC_292_0 (.Y(\u_div/SumTmp[3][2] ), 
	.S0(FE_RN_238_0), 
	.B(FE_RN_239_0), 
	.A(FE_RN_242_0));
   XNOR2X8M FE_RC_291_0 (.Y(FE_RN_237_0), 
	.B(n18), 
	.A(FE_RN_227_0));
   NAND2X4M FE_RC_290_0 (.Y(FE_RN_236_0), 
	.B(FE_RN_230_0), 
	.A(FE_RN_225_0));
   NAND2X4M FE_RC_289_0 (.Y(FE_RN_235_0), 
	.B(\u_div/CryTmp[3][1] ), 
	.A(FE_RN_236_0));
   OAI21X4M FE_RC_288_0 (.Y(\u_div/SumTmp[3][1] ), 
	.B0(FE_RN_235_0), 
	.A1(\u_div/CryTmp[3][1] ), 
	.A0(FE_RN_237_0));
   NOR2BX8M FE_RC_287_0 (.Y(FE_RN_234_0), 
	.B(n17), 
	.AN(FE_RN_230_0));
   NAND2X4M FE_RC_286_0 (.Y(FE_RN_233_0), 
	.B(\u_div/CryTmp[3][1] ), 
	.A(FE_RN_225_0));
   NAND2X4M FE_RC_285_0 (.Y(FE_RN_232_0), 
	.B(FE_RN_234_0), 
	.A(FE_RN_233_0));
   NAND2X4M FE_RC_284_0 (.Y(FE_RN_231_0), 
	.B(\u_div/PartRem[4][2] ), 
	.A(FE_RN_232_0));
   NAND2X8M FE_RC_283_0 (.Y(FE_RN_230_0), 
	.B(n18), 
	.A(FE_RN_227_0));
   CLKNAND2X4M FE_RC_282_0 (.Y(FE_RN_229_0), 
	.B(FE_RN_162_0), 
	.A(FE_RN_189_0));
   NAND2X5M FE_RC_281_0 (.Y(FE_RN_228_0), 
	.B(n21), 
	.A(FE_RN_229_0));
   MXI2X6M FE_RC_280_0 (.Y(FE_RN_227_0), 
	.S0(FE_RN_228_0), 
	.B(FE_RN_191_0), 
	.A(FE_RN_192_0));
   INVX2M FE_RC_279_0 (.Y(FE_RN_226_0), 
	.A(n18));
   NAND2BX8M FE_RC_278_0 (.Y(FE_RN_225_0), 
	.B(FE_RN_226_0), 
	.AN(FE_RN_227_0));
   NAND2X4M FE_RC_277_0 (.Y(FE_RN_224_0), 
	.B(\u_div/CryTmp[3][1] ), 
	.A(FE_RN_225_0));
   NAND2X4M FE_RC_276_0 (.Y(FE_RN_223_0), 
	.B(FE_RN_230_0), 
	.A(FE_RN_224_0));
   NAND2X4M FE_RC_275_0 (.Y(FE_RN_222_0), 
	.B(n17), 
	.A(FE_RN_223_0));
   INVX4M FE_RC_240_0 (.Y(quotient[4]), 
	.A(FE_RN_187_0));
   INVX2M FE_RC_239_0 (.Y(FE_RN_192_0), 
	.A(\u_div/SumTmp[4][0] ));
   INVX2M FE_RC_238_0 (.Y(FE_RN_191_0), 
	.A(a[4]));
   INVX2M FE_RC_237_0 (.Y(FE_RN_190_0), 
	.A(FE_RN_166_0));
   NAND2BX2M FE_RC_236_0 (.Y(FE_RN_189_0), 
	.B(\u_div/CryTmp[4][3] ), 
	.AN(FE_RN_190_0));
   NAND2X2M FE_RC_226_0 (.Y(FE_RN_134_0), 
	.B(FE_RN_135_0), 
	.A(n20));
   INVX2M FE_RC_225_0 (.Y(quotient[5]), 
	.A(FE_RN_164_0));
   NAND2X2M FE_RC_224_0 (.Y(FE_RN_182_0), 
	.B(\u_div/PartRem[6][2] ), 
	.A(FE_RN_164_0));
   INVX2M FE_RC_223_0 (.Y(FE_RN_181_0), 
	.A(FE_RN_165_0));
   CLKNAND2X2M FE_RC_222_0 (.Y(\u_div/PartRem[5][3] ), 
	.B(FE_RN_182_0), 
	.A(FE_RN_181_0));
   INVX2M FE_RC_221_0 (.Y(FE_RN_180_0), 
	.A(\u_div/CryTmp[4][3] ));
   INVX2M FE_RC_220_0 (.Y(FE_RN_179_0), 
	.A(FE_RN_164_0));
   INVX2M FE_RC_219_0 (.Y(FE_RN_178_0), 
	.A(\u_div/PartRem[6][2] ));
   INVX2M FE_RC_218_0 (.Y(FE_RN_177_0), 
	.A(n16));
   OAI22X1M FE_RC_217_0 (.Y(FE_RN_176_0), 
	.B1(\u_div/PartRem[6][2] ), 
	.B0(FE_RN_177_0), 
	.A1(n16), 
	.A0(FE_RN_178_0));
   INVX2M FE_RC_216_0 (.Y(FE_RN_175_0), 
	.A(n16));
   INVX2M FE_RC_215_0 (.Y(FE_RN_174_0), 
	.A(n16));
   OAI2BB2X1M FE_RC_214_0 (.Y(FE_RN_173_0), 
	.B1(FE_RN_174_0), 
	.B0(\u_div/SumTmp[5][2] ), 
	.A1N(\u_div/SumTmp[5][2] ), 
	.A0N(FE_RN_175_0));
   OAI22X1M FE_RC_213_0 (.Y(FE_RN_172_0), 
	.B1(FE_RN_173_0), 
	.B0(FE_RN_164_0), 
	.A1(FE_RN_176_0), 
	.A0(FE_RN_179_0));
   MXI2X2M FE_RC_212_0 (.Y(\u_div/SumTmp[4][3] ), 
	.S0(FE_RN_172_0), 
	.B(FE_RN_180_0), 
	.A(\u_div/CryTmp[4][3] ));
   NAND2BX2M FE_RC_211_0 (.Y(FE_RN_171_0), 
	.B(\u_div/PartRem[6][2] ), 
	.AN(FE_RN_135_0));
   INVX2M FE_RC_210_0 (.Y(FE_RN_170_0), 
	.A(\u_div/PartRem[6][2] ));
   INVX2M FE_RC_209_0 (.Y(FE_RN_169_0), 
	.A(n16));
   OAI21X2M FE_RC_208_0 (.Y(FE_RN_168_0), 
	.B0(FE_RN_169_0), 
	.A1(n20), 
	.A0(FE_RN_170_0));
   NOR2X2M FE_RC_207_0 (.Y(FE_RN_167_0), 
	.B(FE_RN_168_0), 
	.A(FE_RN_165_0));
   NAND2X2M FE_RC_206_0 (.Y(FE_RN_166_0), 
	.B(FE_RN_171_0), 
	.A(FE_RN_167_0));
   NOR2BX2M FE_RC_205_0 (.Y(FE_RN_165_0), 
	.B(FE_RN_164_0), 
	.AN(\u_div/SumTmp[5][2] ));
   NAND2X2M FE_RC_204_0 (.Y(FE_RN_164_0), 
	.B(n20), 
	.A(FE_RN_135_0));
   AND2X2M FE_RC_203_0 (.Y(FE_RN_163_0), 
	.B(\u_div/PartRem[6][2] ), 
	.A(FE_RN_164_0));
   OAI21X2M FE_RC_202_0 (.Y(FE_RN_162_0), 
	.B0(n16), 
	.A1(FE_RN_163_0), 
	.A0(FE_RN_165_0));
   NAND2X5M FE_RC_200_0 (.Y(\u_div/CryTmp[5][3] ), 
	.B(FE_RN_69_0), 
	.A(FE_RN_76_0));
   INVX2M FE_RC_198_0 (.Y(FE_RN_161_0), 
	.A(FE_RN_133_0));
   NAND2X4M FE_RC_197_0 (.Y(FE_RN_160_0), 
	.B(\u_div/PartRem[6][1] ), 
	.A(FE_RN_134_0));
   CLKNAND2X4M FE_RC_196_0 (.Y(\u_div/PartRem[5][2] ), 
	.B(FE_RN_161_0), 
	.A(FE_RN_160_0));
   INVX2M FE_RC_195_0 (.Y(FE_RN_159_0), 
	.A(\u_div/CryTmp[4][2] ));
   INVX2M FE_RC_194_0 (.Y(FE_RN_158_0), 
	.A(\u_div/PartRem[6][1] ));
   INVX2M FE_RC_193_0 (.Y(FE_RN_157_0), 
	.A(n17));
   OAI22X1M FE_RC_192_0 (.Y(FE_RN_156_0), 
	.B1(\u_div/PartRem[6][1] ), 
	.B0(FE_RN_157_0), 
	.A1(n17), 
	.A0(FE_RN_158_0));
   INVX2M FE_RC_191_0 (.Y(FE_RN_155_0), 
	.A(FE_RN_156_0));
   MXI2X2M FE_RC_190_0 (.Y(FE_RN_154_0), 
	.S0(FE_RN_155_0), 
	.B(FE_RN_159_0), 
	.A(\u_div/CryTmp[4][2] ));
   NAND2X3M FE_RC_189_0 (.Y(FE_RN_153_0), 
	.B(FE_RN_134_0), 
	.A(FE_RN_154_0));
   INVX2M FE_RC_188_0 (.Y(FE_RN_152_0), 
	.A(FE_RN_134_0));
   INVX2M FE_RC_187_0 (.Y(FE_RN_151_0), 
	.A(\u_div/CryTmp[4][2] ));
   INVX2M FE_RC_186_0 (.Y(FE_RN_150_0), 
	.A(\u_div/SumTmp[5][1] ));
   INVX2M FE_RC_185_0 (.Y(FE_RN_149_0), 
	.A(n17));
   OAI22X1M FE_RC_184_0 (.Y(FE_RN_148_0), 
	.B1(\u_div/SumTmp[5][1] ), 
	.B0(FE_RN_149_0), 
	.A1(n17), 
	.A0(FE_RN_150_0));
   INVX2M FE_RC_183_0 (.Y(FE_RN_147_0), 
	.A(FE_RN_148_0));
   MXI2X2M FE_RC_182_0 (.Y(FE_RN_146_0), 
	.S0(FE_RN_147_0), 
	.B(FE_RN_151_0), 
	.A(\u_div/CryTmp[4][2] ));
   NAND2X3M FE_RC_181_0 (.Y(FE_RN_145_0), 
	.B(FE_RN_152_0), 
	.A(FE_RN_146_0));
   NAND2X2M FE_RC_180_0 (.Y(\u_div/SumTmp[4][2] ), 
	.B(FE_RN_153_0), 
	.A(FE_RN_145_0));
   INVX2M FE_RC_179_0 (.Y(FE_RN_144_0), 
	.A(FE_RN_135_0));
   INVX2M FE_RC_178_0 (.Y(FE_RN_143_0), 
	.A(\u_div/PartRem[6][1] ));
   INVX2M FE_RC_177_0 (.Y(FE_RN_142_0), 
	.A(\u_div/PartRem[6][1] ));
   INVX2M FE_RC_176_0 (.Y(FE_RN_141_0), 
	.A(n17));
   OAI21X2M FE_RC_175_0 (.Y(FE_RN_140_0), 
	.B0(FE_RN_141_0), 
	.A1(n20), 
	.A0(FE_RN_142_0));
   AOI2B1X2M FE_RC_174_0 (.Y(FE_RN_139_0), 
	.B0(FE_RN_140_0), 
	.A1N(FE_RN_143_0), 
	.A0(FE_RN_144_0));
   OAI2B1X2M FE_RC_173_0 (.Y(FE_RN_138_0), 
	.B0(\u_div/CryTmp[4][2] ), 
	.A1N(FE_RN_139_0), 
	.A0(FE_RN_133_0));
   AND2X4M FE_RC_172_0 (.Y(FE_RN_137_0), 
	.B(\u_div/PartRem[6][1] ), 
	.A(FE_RN_134_0));
   INVX2M FE_RC_171_0 (.Y(FE_RN_136_0), 
	.A(\u_div/SumTmp[5][1] ));
   NAND2X2M FE_RC_170_0 (.Y(FE_RN_135_0), 
	.B(FE_RN_76_0), 
	.A(FE_RN_69_0));
   NOR2X4M FE_RC_168_0 (.Y(FE_RN_133_0), 
	.B(FE_RN_136_0), 
	.A(FE_RN_134_0));
   OAI21X4M FE_RC_167_0 (.Y(FE_RN_132_0), 
	.B0(n17), 
	.A1(FE_RN_133_0), 
	.A0(FE_RN_137_0));
   NAND2X3M FE_RC_166_0 (.Y(\u_div/CryTmp[4][3] ), 
	.B(FE_RN_138_0), 
	.A(FE_RN_132_0));
   NAND2BX2M FE_RC_165_0 (.Y(FE_RN_131_0), 
	.B(\u_div/CryTmp[5][3] ), 
	.AN(FE_RN_110_0));
   OAI2B11X4M FE_RC_164_0 (.Y(\u_div/PartRem[5][1] ), 
	.C0(FE_RN_99_0), 
	.B0(FE_RN_131_0), 
	.A1N(a[5]), 
	.A0(\u_div/CryTmp[5][3] ));
   CLKNAND2X4M FE_RC_163_0 (.Y(FE_RN_130_0), 
	.B(a[5]), 
	.A(FE_RN_116_0));
   INVX2M FE_RC_162_0 (.Y(FE_RN_129_0), 
	.A(a[5]));
   INVX2M FE_RC_161_0 (.Y(FE_RN_128_0), 
	.A(FE_RN_121_0));
   NAND3X3M FE_RC_160_0 (.Y(FE_RN_127_0), 
	.C(FE_RN_99_0), 
	.B(FE_RN_129_0), 
	.A(FE_RN_128_0));
   CLKNAND2X2M FE_RC_159_0 (.Y(FE_RN_126_0), 
	.B(FE_RN_130_0), 
	.A(FE_RN_127_0));
   INVX2M FE_RC_158_0 (.Y(FE_RN_125_0), 
	.A(FE_RN_99_0));
   INVX2M FE_RC_157_0 (.Y(FE_RN_124_0), 
	.A(\u_div/CryTmp[4][1] ));
   INVX2M FE_RC_156_0 (.Y(FE_RN_123_0), 
	.A(n18));
   INVX2M FE_RC_155_0 (.Y(FE_RN_122_0), 
	.A(FE_RN_102_0));
   OAI2BB1X2M FE_RC_154_0 (.Y(FE_RN_121_0), 
	.B0(FE_RN_122_0), 
	.A1N(FE_RN_123_0), 
	.A0N(FE_RN_124_0));
   INVX2M FE_RC_153_0 (.Y(FE_RN_120_0), 
	.A(FE_RN_110_0));
   NOR3X4M FE_RC_152_0 (.Y(FE_RN_119_0), 
	.C(FE_RN_125_0), 
	.B(FE_RN_121_0), 
	.A(FE_RN_120_0));
   NOR2BX8M FE_RC_151_0 (.Y(FE_RN_118_0), 
	.B(FE_RN_110_0), 
	.AN(FE_RN_116_0));
   OAI21X3M FE_RC_150_0 (.Y(FE_RN_117_0), 
	.B0(\u_div/CryTmp[5][3] ), 
	.A1(FE_RN_118_0), 
	.A0(FE_RN_119_0));
   NAND2BX8M FE_RC_149_0 (.Y(FE_RN_116_0), 
	.B(FE_RN_104_0), 
	.AN(FE_RN_102_0));
   NAND2BX8M FE_RC_148_0 (.Y(FE_RN_115_0), 
	.B(FE_RN_116_0), 
	.AN(FE_RN_99_0));
   OAI2B11X2M FE_RC_147_0 (.Y(\u_div/SumTmp[4][1] ), 
	.C0(FE_RN_115_0), 
	.B0(FE_RN_117_0), 
	.A1N(FE_RN_126_0), 
	.A0(\u_div/CryTmp[5][3] ));
   INVX2M FE_RC_146_0 (.Y(FE_RN_114_0), 
	.A(a[5]));
   NOR2BX8M FE_RC_145_0 (.Y(FE_RN_113_0), 
	.B(FE_RN_114_0), 
	.AN(FE_RN_104_0));
   INVX2M FE_RC_144_0 (.Y(FE_RN_112_0), 
	.A(FE_RN_104_0));
   INVX2M FE_RC_143_0 (.Y(FE_RN_111_0), 
	.A(\u_div/SumTmp[5][0] ));
   NAND2BX8M FE_RC_142_0 (.Y(FE_RN_110_0), 
	.B(n20), 
	.AN(FE_RN_111_0));
   INVX2M FE_RC_141_0 (.Y(FE_RN_109_0), 
	.A(FE_RN_110_0));
   NAND2BX2M FE_RC_140_0 (.Y(FE_RN_108_0), 
	.B(FE_RN_109_0), 
	.AN(FE_RN_112_0));
   NAND2BX2M FE_RC_139_0 (.Y(FE_RN_107_0), 
	.B(\u_div/CryTmp[5][3] ), 
	.AN(FE_RN_108_0));
   INVX2M FE_RC_138_0 (.Y(FE_RN_106_0), 
	.A(FE_RN_99_0));
   INVX2M FE_RC_137_0 (.Y(FE_RN_105_0), 
	.A(n18));
   NAND2BX8M FE_RC_136_0 (.Y(FE_RN_104_0), 
	.B(FE_RN_105_0), 
	.AN(\u_div/CryTmp[4][1] ));
   INVX2M FE_RC_135_0 (.Y(FE_RN_103_0), 
	.A(FE_RN_104_0));
   AND2X4M FE_RC_134_0 (.Y(FE_RN_102_0), 
	.B(\u_div/CryTmp[4][1] ), 
	.A(n18));
   AOI2B1X4M FE_RC_133_0 (.Y(FE_RN_101_0), 
	.B0(FE_RN_102_0), 
	.A1N(FE_RN_103_0), 
	.A0(FE_RN_106_0));
   OAI2B11X4M FE_RC_132_0 (.Y(\u_div/CryTmp[4][2] ), 
	.C0(FE_RN_101_0), 
	.B0(FE_RN_107_0), 
	.A1N(FE_RN_113_0), 
	.A0(\u_div/CryTmp[5][3] ));
   NAND2BX8M FE_RC_129_0 (.Y(FE_RN_99_0), 
	.B(a[5]), 
	.AN(n20));
   NAND2X4M FE_RC_109_0 (.Y(FE_RN_41_0), 
	.B(FE_RN_42_0), 
	.A(FE_RN_43_0));
   INVX2M FE_RC_108_0 (.Y(quotient[6]), 
	.A(FE_RN_74_0));
   INVX2M FE_RC_107_0 (.Y(FE_RN_84_0), 
	.A(FE_RN_73_0));
   NAND2X4M FE_RC_106_0 (.Y(FE_RN_83_0), 
	.B(\u_div/PartRem[7][1] ), 
	.A(FE_RN_74_0));
   CLKNAND2X4M FE_RC_105_0 (.Y(\u_div/PartRem[6][2] ), 
	.B(FE_RN_84_0), 
	.A(FE_RN_83_0));
   XOR2X2M FE_RC_104_0 (.Y(FE_RN_82_0), 
	.B(n17), 
	.A(\u_div/SumTmp[6][1] ));
   INVX2M FE_RC_103_0 (.Y(FE_RN_81_0), 
	.A(\u_div/PartRem[7][1] ));
   INVX2M FE_RC_102_0 (.Y(FE_RN_80_0), 
	.A(n17));
   OAI22X1M FE_RC_101_0 (.Y(FE_RN_79_0), 
	.B1(\u_div/PartRem[7][1] ), 
	.B0(FE_RN_80_0), 
	.A1(n17), 
	.A0(FE_RN_81_0));
   MXI2X2M FE_RC_100_0 (.Y(FE_RN_78_0), 
	.S0(FE_RN_74_0), 
	.B(FE_RN_79_0), 
	.A(FE_RN_82_0));
   XNOR2X2M FE_RC_99_0 (.Y(\u_div/SumTmp[5][2] ), 
	.B(\u_div/CryTmp[5][2] ), 
	.A(FE_RN_78_0));
   NAND2X4M FE_RC_98_0 (.Y(FE_RN_77_0), 
	.B(\u_div/PartRem[7][1] ), 
	.A(FE_RN_74_0));
   OAI2B1X4M FE_RC_97_0 (.Y(FE_RN_76_0), 
	.B0(n17), 
	.A1N(FE_RN_77_0), 
	.A0(FE_RN_73_0));
   INVX2M FE_RC_96_0 (.Y(FE_RN_75_0), 
	.A(\u_div/SumTmp[6][1] ));
   NAND2X2M FE_RC_95_0 (.Y(FE_RN_74_0), 
	.B(FE_RN_43_0), 
	.A(FE_RN_42_0));
   NOR2X4M FE_RC_94_0 (.Y(FE_RN_73_0), 
	.B(FE_RN_75_0), 
	.A(FE_RN_74_0));
   INVX2M FE_RC_93_0 (.Y(FE_RN_72_0), 
	.A(\u_div/PartRem[7][1] ));
   AOI2B1X1M FE_RC_92_0 (.Y(FE_RN_71_0), 
	.B0(n17), 
	.A1N(FE_RN_42_0), 
	.A0(\u_div/PartRem[7][1] ));
   OAI21X2M FE_RC_91_0 (.Y(FE_RN_70_0), 
	.B0(FE_RN_71_0), 
	.A1(FE_RN_43_0), 
	.A0(FE_RN_72_0));
   OAI21X3M FE_RC_90_0 (.Y(FE_RN_69_0), 
	.B0(\u_div/CryTmp[5][2] ), 
	.A1(FE_RN_70_0), 
	.A0(FE_RN_73_0));
   MXI2X4M FE_RC_88_0 (.Y(\u_div/PartRem[6][1] ), 
	.S0(FE_RN_41_0), 
	.B(FE_RN_47_0), 
	.A(FE_RN_48_0));
   INVX2M FE_RC_87_0 (.Y(FE_RN_68_0), 
	.A(FE_RN_50_0));
   OAI21X2M FE_RC_86_0 (.Y(FE_RN_67_0), 
	.B0(FE_RN_68_0), 
	.A1(\u_div/CryTmp[5][1] ), 
	.A0(n18));
   NOR2BX8M FE_RC_85_0 (.Y(FE_RN_66_0), 
	.B(FE_RN_50_0), 
	.AN(FE_RN_54_0));
   INVX2M FE_RC_84_0 (.Y(FE_RN_65_0), 
	.A(FE_RN_48_0));
   MXI2X2M FE_RC_83_0 (.Y(FE_RN_64_0), 
	.S0(FE_RN_65_0), 
	.B(FE_RN_66_0), 
	.A(FE_RN_67_0));
   INVX2M FE_RC_82_0 (.Y(FE_RN_63_0), 
	.A(\u_div/CryTmp[5][1] ));
   INVX2M FE_RC_81_0 (.Y(FE_RN_62_0), 
	.A(\u_div/CryTmp[5][1] ));
   NAND2X4M FE_RC_80_0 (.Y(FE_RN_61_0), 
	.B(n18), 
	.A(FE_RN_47_0));
   OAI21X6M FE_RC_79_0 (.Y(FE_RN_60_0), 
	.B0(FE_RN_61_0), 
	.A1(n18), 
	.A0(FE_RN_47_0));
   NAND2X4M FE_RC_78_0 (.Y(FE_RN_59_0), 
	.B(FE_RN_62_0), 
	.A(FE_RN_60_0));
   OAI21X4M FE_RC_77_0 (.Y(FE_RN_58_0), 
	.B0(FE_RN_59_0), 
	.A1(FE_RN_63_0), 
	.A0(FE_RN_60_0));
   CLKNAND2X4M FE_RC_76_0 (.Y(FE_RN_57_0), 
	.B(FE_RN_41_0), 
	.A(FE_RN_58_0));
   OAI2B1X4M FE_RC_75_0 (.Y(\u_div/SumTmp[5][1] ), 
	.B0(FE_RN_57_0), 
	.A1N(FE_RN_64_0), 
	.A0(FE_RN_41_0));
   NOR2BX8M FE_RC_74_0 (.Y(FE_RN_56_0), 
	.B(FE_RN_48_0), 
	.AN(FE_RN_54_0));
   INVX2M FE_RC_73_0 (.Y(FE_RN_55_0), 
	.A(n18));
   NAND2BX8M FE_RC_72_0 (.Y(FE_RN_54_0), 
	.B(FE_RN_55_0), 
	.AN(\u_div/CryTmp[5][1] ));
   NOR2BX8M FE_RC_71_0 (.Y(FE_RN_53_0), 
	.B(FE_RN_47_0), 
	.AN(FE_RN_54_0));
   CLKNAND2X4M FE_RC_70_0 (.Y(FE_RN_52_0), 
	.B(FE_RN_41_0), 
	.A(FE_RN_53_0));
   INVX2M FE_RC_69_0 (.Y(FE_RN_51_0), 
	.A(n18));
   NOR2BX8M FE_RC_68_0 (.Y(FE_RN_50_0), 
	.B(FE_RN_51_0), 
	.AN(\u_div/CryTmp[5][1] ));
   INVX2M FE_RC_67_0 (.Y(FE_RN_49_0), 
	.A(FE_RN_50_0));
   OAI2B11X4M FE_RC_66_0 (.Y(\u_div/CryTmp[5][2] ), 
	.C0(FE_RN_49_0), 
	.B0(FE_RN_52_0), 
	.A1N(FE_RN_56_0), 
	.A0(FE_RN_41_0));
   INVX2M FE_RC_64_0 (.Y(FE_RN_48_0), 
	.A(\u_div/SumTmp[6][0] ));
   INVX2M FE_RC_63_0 (.Y(FE_RN_47_0), 
	.A(a[6]));
   INVX2M FE_RC_62_0 (.Y(FE_RN_46_0), 
	.A(FE_RN_35_0));
   INVX2M FE_RC_61_0 (.Y(FE_RN_45_0), 
	.A(FE_RN_18_0));
   NAND3X3M FE_RC_60_0 (.Y(FE_RN_44_0), 
	.C(FE_RN_38_0), 
	.B(\u_div/SumTmp[7][0] ), 
	.A(FE_RN_45_0));
   NAND3BX2M FE_RC_59_0 (.Y(FE_RN_43_0), 
	.C(FE_RN_34_0), 
	.B(FE_RN_44_0), 
	.AN(FE_RN_46_0));
   NOR2X4M FE_RC_58_0 (.Y(FE_RN_42_0), 
	.B(FE_RN_40_0), 
	.A(FE_RN_39_0));
   INVX2M FE_RC_55_0 (.Y(FE_RN_40_0), 
	.A(n17));
   INVX2M FE_RC_54_0 (.Y(FE_RN_39_0), 
	.A(n20));
   INVX2M FE_RC_53_0 (.Y(FE_RN_38_0), 
	.A(FE_RN_13_0));
   INVX2M FE_RC_52_0 (.Y(FE_RN_37_0), 
	.A(FE_RN_11_0));
   INVX2M FE_RC_51_0 (.Y(FE_RN_36_0), 
	.A(FE_RN_12_0));
   NAND2X3M FE_RC_50_0 (.Y(FE_RN_35_0), 
	.B(FE_RN_37_0), 
	.A(FE_RN_36_0));
   NAND3BX4M FE_RC_49_0 (.Y(FE_RN_34_0), 
	.C(a[7]), 
	.B(FE_RN_18_0), 
	.AN(FE_RN_13_0));
   INVX3M FE_RC_45_0 (.Y(quotient[7]), 
	.A(FE_RN_18_0));
   INVX2M FE_RC_44_0 (.Y(FE_RN_31_0), 
	.A(\u_div/SumTmp[7][0] ));
   NAND2X4M FE_RC_43_0 (.Y(FE_RN_30_0), 
	.B(a[7]), 
	.A(FE_RN_18_0));
   OAI21X4M FE_RC_42_0 (.Y(\u_div/PartRem[7][1] ), 
	.B0(FE_RN_30_0), 
	.A1(FE_RN_31_0), 
	.A0(FE_RN_18_0));
   NOR2X4M FE_RC_41_0 (.Y(FE_RN_29_0), 
	.B(a[7]), 
	.A(FE_RN_25_0));
   AOI21X4M FE_RC_40_0 (.Y(FE_RN_28_0), 
	.B0(FE_RN_29_0), 
	.A1(a[7]), 
	.A0(FE_RN_25_0));
   INVX2M FE_RC_39_0 (.Y(FE_RN_27_0), 
	.A(n18));
   INVX2M FE_RC_38_0 (.Y(FE_RN_26_0), 
	.A(\u_div/CryTmp[6][1] ));
   OAI21X6M FE_RC_37_0 (.Y(FE_RN_25_0), 
	.B0(FE_RN_14_0), 
	.A1(FE_RN_26_0), 
	.A0(FE_RN_27_0));
   NOR2X4M FE_RC_36_0 (.Y(FE_RN_24_0), 
	.B(\u_div/SumTmp[7][0] ), 
	.A(FE_RN_25_0));
   AOI21X4M FE_RC_35_0 (.Y(FE_RN_23_0), 
	.B0(FE_RN_24_0), 
	.A1(\u_div/SumTmp[7][0] ), 
	.A0(FE_RN_25_0));
   INVX2M FE_RC_34_0 (.Y(FE_RN_22_0), 
	.A(FE_RN_18_0));
   MXI2X4M FE_RC_33_0 (.Y(\u_div/SumTmp[6][1] ), 
	.S0(FE_RN_22_0), 
	.B(FE_RN_23_0), 
	.A(FE_RN_28_0));
   INVX2M FE_RC_31_0 (.Y(FE_RN_20_0), 
	.A(FE_RN_4_0));
   NOR2X3M FE_RC_30_0 (.Y(FE_RN_19_0), 
	.B(FE_RN_5_0), 
	.A(FE_RN_3_0));
   NAND4X6M FE_RC_29_0 (.Y(FE_RN_18_0), 
	.D(FE_RN_20_0), 
	.C(\u_div/CryTmp[7][1] ), 
	.B(n21), 
	.A(FE_RN_19_0));
   INVX2M FE_RC_27_0 (.Y(FE_RN_16_0), 
	.A(\u_div/CryTmp[6][1] ));
   INVX2M FE_RC_26_0 (.Y(FE_RN_15_0), 
	.A(n18));
   NAND2X4M FE_RC_25_0 (.Y(FE_RN_14_0), 
	.B(FE_RN_16_0), 
	.A(FE_RN_15_0));
   INVX2M FE_RC_24_0 (.Y(FE_RN_13_0), 
	.A(FE_RN_14_0));
   INVX2M FE_RC_23_0 (.Y(FE_RN_12_0), 
	.A(\u_div/CryTmp[6][1] ));
   INVX2M FE_RC_22_0 (.Y(FE_RN_11_0), 
	.A(n18));
   AND2X8M FE_RC_13_0 (.Y(n20), 
	.B(n16), 
	.A(n21));
   INVX2M FE_RC_12_0 (.Y(FE_RN_5_0), 
	.A(n17));
   INVX2M FE_RC_11_0 (.Y(FE_RN_4_0), 
	.A(n18));
   INVX2M FE_RC_10_0 (.Y(FE_RN_3_0), 
	.A(n16));
   NOR2X12M FE_RC_7_0 (.Y(n22), 
	.B(b[7]), 
	.A(b[6]));
   NOR2X12M FE_RC_6_0 (.Y(FE_RN_1_0), 
	.B(b[7]), 
	.A(b[6]));
   AND3X6M FE_RC_5_0 (.Y(n21), 
	.C(FE_RN_0_0), 
	.B(n15), 
	.A(FE_RN_1_0));
   INVX10M FE_RC_3_0 (.Y(n14), 
	.A(b[5]));
   INVX2M FE_RC_2_0 (.Y(FE_RN_0_0), 
	.A(b[5]));
   INVX8M FE_RC_0_0 (.Y(n15), 
	.A(b[4]));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_5  (.CO(\u_div/CryTmp[0][6] ), 
	.CI(\u_div/CryTmp[0][5] ), 
	.B(n14), 
	.A(\u_div/PartRem[1][5] ));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_6  (.CO(\u_div/CryTmp[0][7] ), 
	.CI(\u_div/CryTmp[0][6] ), 
	.B(n173), 
	.A(\u_div/PartRem[1][6] ));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_3  (.CO(\u_div/CryTmp[0][4] ), 
	.CI(\u_div/CryTmp[0][3] ), 
	.B(n16), 
	.A(\u_div/PartRem[1][3] ));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_4  (.CO(\u_div/CryTmp[0][5] ), 
	.CI(\u_div/CryTmp[0][4] ), 
	.B(n15), 
	.A(\u_div/PartRem[1][4] ));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_1  (.CO(\u_div/CryTmp[0][2] ), 
	.CI(\u_div/CryTmp[0][1] ), 
	.B(n18), 
	.A(\u_div/PartRem[1][1] ));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_2  (.CO(\u_div/CryTmp[0][3] ), 
	.CI(\u_div/CryTmp[0][2] ), 
	.B(n17), 
	.A(\u_div/PartRem[1][2] ));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_7  (.CO(quotient[0]), 
	.CI(\u_div/CryTmp[0][7] ), 
	.B(n12), 
	.A(\u_div/PartRem[1][7] ));
   INVX12M U1 (.Y(n19), 
	.A(b[0]));
   XNOR2X2M U2 (.Y(\u_div/SumTmp[7][0] ), 
	.B(a[7]), 
	.A(n19));
   XNOR2X2M U3 (.Y(\u_div/SumTmp[6][0] ), 
	.B(a[6]), 
	.A(n19));
   XNOR2X2M U4 (.Y(\u_div/SumTmp[5][0] ), 
	.B(a[5]), 
	.A(n19));
   XNOR2X2M U5 (.Y(\u_div/SumTmp[4][0] ), 
	.B(a[4]), 
	.A(n19));
   XNOR2X2M U6 (.Y(\u_div/SumTmp[3][0] ), 
	.B(a[3]), 
	.A(n19));
   XNOR2X2M U7 (.Y(\u_div/SumTmp[2][0] ), 
	.B(a[2]), 
	.A(n19));
   XNOR2X2M U8 (.Y(\u_div/SumTmp[1][0] ), 
	.B(a[1]), 
	.A(n19));
   OR2X2M U9 (.Y(\u_div/CryTmp[7][1] ), 
	.B(a[7]), 
	.A(n19));
   NAND2X2M U10 (.Y(\u_div/CryTmp[0][1] ), 
	.B(n11), 
	.A(n7));
   NAND2X2M U11 (.Y(\u_div/CryTmp[5][1] ), 
	.B(n4), 
	.A(n3));
   CLKINVX2M U12 (.Y(n4), 
	.A(a[5]));
   CLKINVX2M U13 (.Y(n3), 
	.A(n19));
   NAND2X2M U14 (.Y(\u_div/CryTmp[4][1] ), 
	.B(n6), 
	.A(n5));
   CLKINVX2M U15 (.Y(n6), 
	.A(a[4]));
   CLKINVX2M U16 (.Y(n5), 
	.A(n19));
   NAND2X2M U17 (.Y(\u_div/CryTmp[3][1] ), 
	.B(n8), 
	.A(n7));
   CLKINVX2M U18 (.Y(n8), 
	.A(a[3]));
   INVX2M U19 (.Y(n7), 
	.A(n19));
   NAND2X2M U20 (.Y(\u_div/CryTmp[2][1] ), 
	.B(n9), 
	.A(n7));
   INVX2M U21 (.Y(n9), 
	.A(a[2]));
   NAND2X2M U22 (.Y(\u_div/CryTmp[1][1] ), 
	.B(n10), 
	.A(n7));
   INVX2M U23 (.Y(n10), 
	.A(a[1]));
   NAND2X2M U24 (.Y(\u_div/CryTmp[6][1] ), 
	.B(n2), 
	.A(n1));
   CLKINVX2M U25 (.Y(n2), 
	.A(a[6]));
   CLKINVX2M U26 (.Y(n1), 
	.A(n19));
   INVX2M U27 (.Y(n11), 
	.A(a[0]));
   INVX12M U28 (.Y(n18), 
	.A(b[1]));
   INVX12M U29 (.Y(n17), 
	.A(b[2]));
   INVX8M U30 (.Y(n16), 
	.A(b[3]));
   INVX2M U34 (.Y(n12), 
	.A(b[7]));
   CLKMX2X2M U35 (.Y(\u_div/PartRem[1][7] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][6] ), 
	.A(\u_div/PartRem[2][6] ));
   CLKMX2X2M U36 (.Y(\u_div/PartRem[2][6] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][5] ), 
	.A(\u_div/PartRem[3][5] ));
   CLKMX2X2M U37 (.Y(\u_div/PartRem[3][5] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][4] ), 
	.A(\u_div/PartRem[4][4] ));
   CLKMX2X2M U38 (.Y(\u_div/PartRem[4][4] ), 
	.S0(quotient[4]), 
	.B(\u_div/SumTmp[4][3] ), 
	.A(\u_div/PartRem[5][3] ));
   CLKMX2X2M U42 (.Y(\u_div/PartRem[1][6] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][5] ), 
	.A(\u_div/PartRem[2][5] ));
   CLKMX2X2M U43 (.Y(\u_div/PartRem[2][5] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][4] ), 
	.A(\u_div/PartRem[3][4] ));
   CLKMX2X2M U44 (.Y(\u_div/PartRem[3][4] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][3] ), 
	.A(\u_div/PartRem[4][3] ));
   CLKMX2X2M U45 (.Y(\u_div/PartRem[4][3] ), 
	.S0(quotient[4]), 
	.B(\u_div/SumTmp[4][2] ), 
	.A(\u_div/PartRem[5][2] ));
   CLKMX2X2M U48 (.Y(\u_div/PartRem[1][5] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][4] ), 
	.A(\u_div/PartRem[2][4] ));
   CLKMX2X2M U49 (.Y(\u_div/PartRem[2][4] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][3] ), 
	.A(\u_div/PartRem[3][3] ));
   CLKMX2X2M U50 (.Y(\u_div/PartRem[3][3] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][2] ), 
	.A(\u_div/PartRem[4][2] ));
   CLKMX2X2M U51 (.Y(\u_div/PartRem[4][2] ), 
	.S0(quotient[4]), 
	.B(\u_div/SumTmp[4][1] ), 
	.A(\u_div/PartRem[5][1] ));
   CLKMX2X2M U53 (.Y(\u_div/PartRem[1][4] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][3] ), 
	.A(\u_div/PartRem[2][3] ));
   CLKMX2X2M U54 (.Y(\u_div/PartRem[2][3] ), 
	.S0(quotient[2]), 
	.B(\u_div/SumTmp[2][2] ), 
	.A(\u_div/PartRem[3][2] ));
   CLKMX2X2M U55 (.Y(\u_div/PartRem[3][2] ), 
	.S0(quotient[3]), 
	.B(\u_div/SumTmp[3][1] ), 
	.A(\u_div/PartRem[4][1] ));
   CLKMX2X2M U57 (.Y(\u_div/PartRem[1][3] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][2] ), 
	.A(\u_div/PartRem[2][2] ));
   CLKMX2X2M U60 (.Y(\u_div/PartRem[1][2] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][1] ), 
	.A(\u_div/PartRem[2][1] ));
   MX2X2M U62 (.Y(\u_div/PartRem[1][1] ), 
	.S0(quotient[1]), 
	.B(\u_div/SumTmp[1][0] ), 
	.A(a[1]));
endmodule

module ALU_00000008_00000004_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n170, 
	n173, 
	n172, 
	n195, 
	n171);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n170;
   input n173;
   input n172;
   input n195;
   input n171;

   // Internal wires
   wire n1;
   wire n2;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [9:0] carry;

   ADDFX2M U2_7 (.S(DIFF[7]), 
	.CO(carry[8]), 
	.CI(carry[7]), 
	.B(n2), 
	.A(A[7]));
   ADDFX2M U2_1 (.S(DIFF[1]), 
	.CO(carry[2]), 
	.CI(carry[1]), 
	.B(n8), 
	.A(A[1]));
   ADDFX2M U2_6 (.S(DIFF[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(n173), 
	.A(A[6]));
   ADDFX2M U2_5 (.S(DIFF[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(n4), 
	.A(A[5]));
   ADDFX2M U2_4 (.S(DIFF[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(n5), 
	.A(A[4]));
   ADDFX2M U2_3 (.S(DIFF[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(n6), 
	.A(A[3]));
   ADDFX2M U2_2 (.S(DIFF[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(n7), 
	.A(A[2]));
   XNOR2X2M U1 (.Y(DIFF[0]), 
	.B(A[0]), 
	.A(n9));
   INVX2M U2 (.Y(n9), 
	.A(B[0]));
   INVX2M U3 (.Y(n7), 
	.A(B[2]));
   INVX2M U4 (.Y(n6), 
	.A(B[3]));
   INVX2M U5 (.Y(n5), 
	.A(B[4]));
   INVX2M U6 (.Y(n4), 
	.A(B[5]));
   INVX2M U8 (.Y(n8), 
	.A(B[1]));
   NAND2X2M U9 (.Y(carry[1]), 
	.B(n1), 
	.A(B[0]));
   INVX2M U10 (.Y(n1), 
	.A(A[0]));
   INVX2M U11 (.Y(n2), 
	.A(B[7]));
   CLKINVX1M U12 (.Y(DIFF[8]), 
	.A(carry[8]));
endmodule

module ALU_00000008_00000004_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   ADDFX2M U1_7 (.S(SUM[7]), 
	.CO(SUM[8]), 
	.CI(carry[7]), 
	.B(B[7]), 
	.A(A[7]));
   ADDFX2M U1_1 (.S(SUM[1]), 
	.CO(carry[2]), 
	.CI(n1), 
	.B(B[1]), 
	.A(A[1]));
   ADDFX2M U1_6 (.S(SUM[6]), 
	.CO(carry[7]), 
	.CI(carry[6]), 
	.B(B[6]), 
	.A(A[6]));
   ADDFX2M U1_5 (.S(SUM[5]), 
	.CO(carry[6]), 
	.CI(carry[5]), 
	.B(B[5]), 
	.A(A[5]));
   ADDFX2M U1_4 (.S(SUM[4]), 
	.CO(carry[5]), 
	.CI(carry[4]), 
	.B(B[4]), 
	.A(A[4]));
   ADDFX2M U1_3 (.S(SUM[3]), 
	.CO(carry[4]), 
	.CI(carry[3]), 
	.B(B[3]), 
	.A(A[3]));
   ADDFX2M U1_2 (.S(SUM[2]), 
	.CO(carry[3]), 
	.CI(carry[2]), 
	.B(B[2]), 
	.A(A[2]));
   AND2X2M U1 (.Y(n1), 
	.B(A[0]), 
	.A(B[0]));
   CLKXOR2X2M U2 (.Y(SUM[0]), 
	.B(A[0]), 
	.A(B[0]));
endmodule

module ALU_00000008_00000004_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;

   AOI21BX2M U2 (.Y(n1), 
	.B0N(n19), 
	.A1(A[12]), 
	.A0(n18));
   NAND2X2M U3 (.Y(n15), 
	.B(B[7]), 
	.A(A[7]));
   INVX2M U4 (.Y(n9), 
	.A(A[6]));
   XNOR2X2M U5 (.Y(SUM[13]), 
	.B(n1), 
	.A(B[13]));
   XNOR2X2M U6 (.Y(SUM[7]), 
	.B(n8), 
	.A(A[7]));
   INVX2M U7 (.Y(n8), 
	.A(B[7]));
   INVX2M U8 (.Y(SUM[6]), 
	.A(n9));
   BUFX2M U9 (.Y(SUM[0]), 
	.A(A[0]));
   BUFX2M U10 (.Y(SUM[1]), 
	.A(A[1]));
   BUFX2M U11 (.Y(SUM[2]), 
	.A(A[2]));
   BUFX2M U12 (.Y(SUM[3]), 
	.A(A[3]));
   BUFX2M U13 (.Y(SUM[4]), 
	.A(A[4]));
   BUFX2M U14 (.Y(SUM[5]), 
	.A(A[5]));
   XNOR2X1M U15 (.Y(SUM[9]), 
	.B(n11), 
	.A(n10));
   NOR2X1M U16 (.Y(n11), 
	.B(n13), 
	.A(n12));
   CLKXOR2X2M U17 (.Y(SUM[8]), 
	.B(n15), 
	.A(n14));
   NAND2BX1M U18 (.Y(n14), 
	.B(n17), 
	.AN(n16));
   OAI21X1M U19 (.Y(n19), 
	.B0(B[12]), 
	.A1(n18), 
	.A0(A[12]));
   XOR3XLM U20 (.Y(SUM[12]), 
	.C(n18), 
	.B(A[12]), 
	.A(B[12]));
   OAI21BX1M U21 (.Y(n18), 
	.B0N(n22), 
	.A1(n21), 
	.A0(n20));
   XNOR2X1M U22 (.Y(SUM[11]), 
	.B(n23), 
	.A(n21));
   NOR2X1M U23 (.Y(n23), 
	.B(n20), 
	.A(n22));
   NOR2X1M U24 (.Y(n20), 
	.B(A[11]), 
	.A(B[11]));
   AND2X1M U25 (.Y(n22), 
	.B(A[11]), 
	.A(B[11]));
   OA21X1M U26 (.Y(n21), 
	.B0(n26), 
	.A1(n25), 
	.A0(n24));
   CLKXOR2X2M U27 (.Y(SUM[10]), 
	.B(n25), 
	.A(n27));
   AOI2BB1X1M U28 (.Y(n25), 
	.B0(n12), 
	.A1N(n13), 
	.A0N(n10));
   AND2X1M U29 (.Y(n12), 
	.B(A[9]), 
	.A(B[9]));
   NOR2X1M U30 (.Y(n13), 
	.B(A[9]), 
	.A(B[9]));
   OA21X1M U31 (.Y(n10), 
	.B0(n17), 
	.A1(n16), 
	.A0(n15));
   CLKNAND2X2M U32 (.Y(n17), 
	.B(A[8]), 
	.A(B[8]));
   NOR2X1M U33 (.Y(n16), 
	.B(A[8]), 
	.A(B[8]));
   NAND2BX1M U34 (.Y(n27), 
	.B(n26), 
	.AN(n24));
   CLKNAND2X2M U35 (.Y(n26), 
	.B(A[10]), 
	.A(B[10]));
   NOR2X1M U36 (.Y(n24), 
	.B(A[10]), 
	.A(B[10]));
endmodule

module ALU_00000008_00000004_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n170, 
	n172, 
	n189, 
	n190, 
	n175, 
	n195, 
	n171, 
	n191, 
	n192, 
	n193, 
	n194, 
	n173);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n170;
   input n172;
   input n189;
   input n190;
   input n175;
   input n195;
   input n171;
   input n191;
   input n192;
   input n193;
   input n194;
   input n173;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n30;
   wire n31;
   wire n32;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;

   ADDFX2M S1_2_0 (.S(\A1[0] ), 
	.CO(\CARRYB[2][0] ), 
	.CI(\SUMB[1][1] ), 
	.B(n7), 
	.A(\ab[2][0] ));
   ADDFX2M S3_6_6 (.S(\SUMB[6][6] ), 
	.CO(\CARRYB[6][6] ), 
	.CI(\ab[5][7] ), 
	.B(\CARRYB[5][6] ), 
	.A(\ab[6][6] ));
   ADDFX2M S3_5_6 (.S(\SUMB[5][6] ), 
	.CO(\CARRYB[5][6] ), 
	.CI(\ab[4][7] ), 
	.B(\CARRYB[4][6] ), 
	.A(\ab[5][6] ));
   ADDFX2M S5_6 (.S(\SUMB[7][6] ), 
	.CO(\CARRYB[7][6] ), 
	.CI(\ab[6][7] ), 
	.B(\CARRYB[6][6] ), 
	.A(\ab[7][6] ));
   ADDFX2M S4_5 (.S(\SUMB[7][5] ), 
	.CO(\CARRYB[7][5] ), 
	.CI(\SUMB[6][6] ), 
	.B(\CARRYB[6][5] ), 
	.A(\ab[7][5] ));
   ADDFX2M S1_6_0 (.S(\A1[4] ), 
	.CO(\CARRYB[6][0] ), 
	.CI(\SUMB[5][1] ), 
	.B(\CARRYB[5][0] ), 
	.A(\ab[6][0] ));
   ADDFX2M S2_6_2 (.S(\SUMB[6][2] ), 
	.CO(\CARRYB[6][2] ), 
	.CI(\SUMB[5][3] ), 
	.B(\CARRYB[5][2] ), 
	.A(\ab[6][2] ));
   ADDFX2M S2_6_1 (.S(\SUMB[6][1] ), 
	.CO(\CARRYB[6][1] ), 
	.CI(\SUMB[5][2] ), 
	.B(\CARRYB[5][1] ), 
	.A(\ab[6][1] ));
   ADDFX2M S1_5_0 (.S(\A1[3] ), 
	.CO(\CARRYB[5][0] ), 
	.CI(\SUMB[4][1] ), 
	.B(\CARRYB[4][0] ), 
	.A(\ab[5][0] ));
   ADDFX2M S2_5_3 (.S(\SUMB[5][3] ), 
	.CO(\CARRYB[5][3] ), 
	.CI(\SUMB[4][4] ), 
	.B(\CARRYB[4][3] ), 
	.A(\ab[5][3] ));
   ADDFX2M S2_5_2 (.S(\SUMB[5][2] ), 
	.CO(\CARRYB[5][2] ), 
	.CI(\SUMB[4][3] ), 
	.B(\CARRYB[4][2] ), 
	.A(\ab[5][2] ));
   ADDFX2M S2_5_1 (.S(\SUMB[5][1] ), 
	.CO(\CARRYB[5][1] ), 
	.CI(\SUMB[4][2] ), 
	.B(\CARRYB[4][1] ), 
	.A(\ab[5][1] ));
   ADDFX2M S1_4_0 (.S(\A1[2] ), 
	.CO(\CARRYB[4][0] ), 
	.CI(\SUMB[3][1] ), 
	.B(\CARRYB[3][0] ), 
	.A(\ab[4][0] ));
   ADDFX2M S2_4_4 (.S(\SUMB[4][4] ), 
	.CO(\CARRYB[4][4] ), 
	.CI(\SUMB[3][5] ), 
	.B(\CARRYB[3][4] ), 
	.A(\ab[4][4] ));
   ADDFX2M S2_4_3 (.S(\SUMB[4][3] ), 
	.CO(\CARRYB[4][3] ), 
	.CI(\SUMB[3][4] ), 
	.B(\CARRYB[3][3] ), 
	.A(\ab[4][3] ));
   ADDFX2M S2_4_2 (.S(\SUMB[4][2] ), 
	.CO(\CARRYB[4][2] ), 
	.CI(\SUMB[3][3] ), 
	.B(\CARRYB[3][2] ), 
	.A(\ab[4][2] ));
   ADDFX2M S2_4_1 (.S(\SUMB[4][1] ), 
	.CO(\CARRYB[4][1] ), 
	.CI(\SUMB[3][2] ), 
	.B(\CARRYB[3][1] ), 
	.A(\ab[4][1] ));
   ADDFX2M S1_3_0 (.S(\A1[1] ), 
	.CO(\CARRYB[3][0] ), 
	.CI(\SUMB[2][1] ), 
	.B(\CARRYB[2][0] ), 
	.A(\ab[3][0] ));
   ADDFX2M S2_3_4 (.S(\SUMB[3][4] ), 
	.CO(\CARRYB[3][4] ), 
	.CI(\SUMB[2][5] ), 
	.B(\CARRYB[2][4] ), 
	.A(\ab[3][4] ));
   ADDFX2M S2_3_2 (.S(\SUMB[3][2] ), 
	.CO(\CARRYB[3][2] ), 
	.CI(\SUMB[2][3] ), 
	.B(\CARRYB[2][2] ), 
	.A(\ab[3][2] ));
   ADDFX2M S2_3_1 (.S(\SUMB[3][1] ), 
	.CO(\CARRYB[3][1] ), 
	.CI(\SUMB[2][2] ), 
	.B(\CARRYB[2][1] ), 
	.A(\ab[3][1] ));
   ADDFX2M S2_3_5 (.S(\SUMB[3][5] ), 
	.CO(\CARRYB[3][5] ), 
	.CI(\SUMB[2][6] ), 
	.B(\CARRYB[2][5] ), 
	.A(\ab[3][5] ));
   ADDFX2M S2_2_2 (.S(\SUMB[2][2] ), 
	.CO(\CARRYB[2][2] ), 
	.CI(\SUMB[1][3] ), 
	.B(n6), 
	.A(\ab[2][2] ));
   ADDFX2M S2_2_1 (.S(\SUMB[2][1] ), 
	.CO(\CARRYB[2][1] ), 
	.CI(\SUMB[1][2] ), 
	.B(n5), 
	.A(\ab[2][1] ));
   ADDFX2M S2_6_4 (.S(\SUMB[6][4] ), 
	.CO(\CARRYB[6][4] ), 
	.CI(\SUMB[5][5] ), 
	.B(\CARRYB[5][4] ), 
	.A(\ab[6][4] ));
   ADDFX2M S2_6_3 (.S(\SUMB[6][3] ), 
	.CO(\CARRYB[6][3] ), 
	.CI(\SUMB[5][4] ), 
	.B(\CARRYB[5][3] ), 
	.A(\ab[6][3] ));
   ADDFX2M S2_6_5 (.S(\SUMB[6][5] ), 
	.CO(\CARRYB[6][5] ), 
	.CI(\SUMB[5][6] ), 
	.B(\CARRYB[5][5] ), 
	.A(\ab[6][5] ));
   ADDFX2M S2_5_4 (.S(\SUMB[5][4] ), 
	.CO(\CARRYB[5][4] ), 
	.CI(\SUMB[4][5] ), 
	.B(\CARRYB[4][4] ), 
	.A(\ab[5][4] ));
   ADDFX2M S2_5_5 (.S(\SUMB[5][5] ), 
	.CO(\CARRYB[5][5] ), 
	.CI(\SUMB[4][6] ), 
	.B(\CARRYB[4][5] ), 
	.A(\ab[5][5] ));
   ADDFX2M S3_4_6 (.S(\SUMB[4][6] ), 
	.CO(\CARRYB[4][6] ), 
	.CI(\ab[3][7] ), 
	.B(\CARRYB[3][6] ), 
	.A(\ab[4][6] ));
   ADDFX2M S2_4_5 (.S(\SUMB[4][5] ), 
	.CO(\CARRYB[4][5] ), 
	.CI(\SUMB[3][6] ), 
	.B(\CARRYB[3][5] ), 
	.A(\ab[4][5] ));
   ADDFX2M S2_3_3 (.S(\SUMB[3][3] ), 
	.CO(\CARRYB[3][3] ), 
	.CI(\SUMB[2][4] ), 
	.B(\CARRYB[2][3] ), 
	.A(\ab[3][3] ));
   ADDFX2M S3_3_6 (.S(\SUMB[3][6] ), 
	.CO(\CARRYB[3][6] ), 
	.CI(\ab[2][7] ), 
	.B(\CARRYB[2][6] ), 
	.A(\ab[3][6] ));
   ADDFX2M S2_2_3 (.S(\SUMB[2][3] ), 
	.CO(\CARRYB[2][3] ), 
	.CI(\SUMB[1][4] ), 
	.B(n4), 
	.A(\ab[2][3] ));
   ADDFX2M S3_2_6 (.S(\SUMB[2][6] ), 
	.CO(\CARRYB[2][6] ), 
	.CI(\ab[1][7] ), 
	.B(n9), 
	.A(\ab[2][6] ));
   ADDFX2M S2_2_5 (.S(\SUMB[2][5] ), 
	.CO(\CARRYB[2][5] ), 
	.CI(\SUMB[1][6] ), 
	.B(n8), 
	.A(\ab[2][5] ));
   ADDFX2M S4_0 (.S(\SUMB[7][0] ), 
	.CO(\CARRYB[7][0] ), 
	.CI(\SUMB[6][1] ), 
	.B(\CARRYB[6][0] ), 
	.A(\ab[7][0] ));
   ADDFX2M S4_4 (.S(\SUMB[7][4] ), 
	.CO(\CARRYB[7][4] ), 
	.CI(\SUMB[6][5] ), 
	.B(\CARRYB[6][4] ), 
	.A(\ab[7][4] ));
   ADDFX2M S4_3 (.S(\SUMB[7][3] ), 
	.CO(\CARRYB[7][3] ), 
	.CI(\SUMB[6][4] ), 
	.B(\CARRYB[6][3] ), 
	.A(\ab[7][3] ));
   ADDFX2M S4_2 (.S(\SUMB[7][2] ), 
	.CO(\CARRYB[7][2] ), 
	.CI(\SUMB[6][3] ), 
	.B(\CARRYB[6][2] ), 
	.A(\ab[7][2] ));
   ADDFX2M S4_1 (.S(\SUMB[7][1] ), 
	.CO(\CARRYB[7][1] ), 
	.CI(\SUMB[6][2] ), 
	.B(\CARRYB[6][1] ), 
	.A(\ab[7][1] ));
   ADDFX2M S2_2_4 (.S(\SUMB[2][4] ), 
	.CO(\CARRYB[2][4] ), 
	.CI(\SUMB[1][5] ), 
	.B(n3), 
	.A(\ab[2][4] ));
   AND2X2M U2 (.Y(n3), 
	.B(\ab[1][4] ), 
	.A(\ab[0][5] ));
   AND2X2M U3 (.Y(n4), 
	.B(\ab[1][3] ), 
	.A(\ab[0][4] ));
   AND2X2M U4 (.Y(n5), 
	.B(\ab[1][1] ), 
	.A(\ab[0][2] ));
   AND2X2M U5 (.Y(n6), 
	.B(\ab[1][2] ), 
	.A(\ab[0][3] ));
   AND2X2M U6 (.Y(n7), 
	.B(\ab[1][0] ), 
	.A(\ab[0][1] ));
   AND2X2M U7 (.Y(n8), 
	.B(\ab[1][5] ), 
	.A(\ab[0][6] ));
   AND2X2M U8 (.Y(n9), 
	.B(\ab[1][6] ), 
	.A(\ab[0][7] ));
   AND2X2M U9 (.Y(n10), 
	.B(\ab[7][7] ), 
	.A(\CARRYB[7][6] ));
   CLKXOR2X2M U10 (.Y(\A1[7] ), 
	.B(\SUMB[7][2] ), 
	.A(\CARRYB[7][1] ));
   CLKXOR2X2M U11 (.Y(\A1[8] ), 
	.B(\SUMB[7][3] ), 
	.A(\CARRYB[7][2] ));
   CLKXOR2X2M U12 (.Y(\A1[9] ), 
	.B(\SUMB[7][4] ), 
	.A(\CARRYB[7][3] ));
   INVX2M U13 (.Y(n23), 
	.A(\ab[0][7] ));
   INVX2M U14 (.Y(n19), 
	.A(\ab[0][3] ));
   INVX2M U15 (.Y(n20), 
	.A(\ab[0][4] ));
   INVX2M U16 (.Y(n21), 
	.A(\ab[0][5] ));
   INVX2M U17 (.Y(n22), 
	.A(\ab[0][6] ));
   AND2X2M U18 (.Y(n11), 
	.B(\SUMB[7][1] ), 
	.A(\CARRYB[7][0] ));
   AND2X2M U19 (.Y(n12), 
	.B(\SUMB[7][2] ), 
	.A(\CARRYB[7][1] ));
   AND2X2M U20 (.Y(n13), 
	.B(\SUMB[7][3] ), 
	.A(\CARRYB[7][2] ));
   CLKXOR2X2M U21 (.Y(\A1[10] ), 
	.B(\SUMB[7][5] ), 
	.A(\CARRYB[7][4] ));
   CLKXOR2X2M U22 (.Y(\A1[11] ), 
	.B(\SUMB[7][6] ), 
	.A(\CARRYB[7][5] ));
   INVX2M U23 (.Y(n18), 
	.A(\ab[0][2] ));
   AND2X2M U24 (.Y(n14), 
	.B(\SUMB[7][4] ), 
	.A(\CARRYB[7][3] ));
   AND2X2M U25 (.Y(n15), 
	.B(\SUMB[7][6] ), 
	.A(\CARRYB[7][5] ));
   AND2X2M U26 (.Y(n16), 
	.B(\SUMB[7][5] ), 
	.A(\CARRYB[7][4] ));
   CLKXOR2X2M U27 (.Y(\A1[12] ), 
	.B(\ab[7][7] ), 
	.A(\CARRYB[7][6] ));
   XNOR2X2M U28 (.Y(\A1[6] ), 
	.B(n17), 
	.A(\CARRYB[7][0] ));
   INVX2M U29 (.Y(n17), 
	.A(\SUMB[7][1] ));
   CLKXOR2X2M U30 (.Y(PRODUCT[1]), 
	.B(\ab[0][1] ), 
	.A(\ab[1][0] ));
   XNOR2X2M U31 (.Y(\SUMB[1][5] ), 
	.B(n22), 
	.A(\ab[1][5] ));
   XNOR2X2M U32 (.Y(\SUMB[1][6] ), 
	.B(n23), 
	.A(\ab[1][6] ));
   XNOR2X2M U33 (.Y(\SUMB[1][4] ), 
	.B(n21), 
	.A(\ab[1][4] ));
   XNOR2X2M U34 (.Y(\SUMB[1][2] ), 
	.B(n19), 
	.A(\ab[1][2] ));
   XNOR2X2M U35 (.Y(\SUMB[1][3] ), 
	.B(n20), 
	.A(\ab[1][3] ));
   INVX2M U36 (.Y(n30), 
	.A(A[1]));
   INVX2M U37 (.Y(n31), 
	.A(A[0]));
   XNOR2X2M U39 (.Y(\SUMB[1][1] ), 
	.B(n18), 
	.A(\ab[1][1] ));
   INVX2M U46 (.Y(n37), 
	.A(B[2]));
   INVX2M U47 (.Y(n36), 
	.A(B[3]));
   INVX2M U48 (.Y(n32), 
	.A(B[7]));
   INVX2M U49 (.Y(n35), 
	.A(B[4]));
   INVX2M U50 (.Y(n34), 
	.A(B[5]));
   INVX2M U51 (.Y(n39), 
	.A(B[0]));
   INVX2M U52 (.Y(n38), 
	.A(B[1]));
   NOR2X1M U54 (.Y(\ab[7][7] ), 
	.B(n32), 
	.A(n189));
   NOR2X1M U55 (.Y(\ab[7][6] ), 
	.B(n173), 
	.A(n189));
   NOR2X1M U56 (.Y(\ab[7][5] ), 
	.B(n34), 
	.A(n189));
   NOR2X1M U57 (.Y(\ab[7][4] ), 
	.B(n35), 
	.A(n189));
   NOR2X1M U58 (.Y(\ab[7][3] ), 
	.B(n36), 
	.A(n189));
   NOR2X1M U59 (.Y(\ab[7][2] ), 
	.B(n37), 
	.A(n189));
   NOR2X1M U60 (.Y(\ab[7][1] ), 
	.B(n38), 
	.A(n189));
   NOR2X1M U61 (.Y(\ab[7][0] ), 
	.B(n39), 
	.A(n189));
   NOR2X1M U62 (.Y(\ab[6][7] ), 
	.B(n190), 
	.A(n32));
   NOR2X1M U63 (.Y(\ab[6][6] ), 
	.B(n190), 
	.A(n173));
   NOR2X1M U64 (.Y(\ab[6][5] ), 
	.B(n190), 
	.A(n34));
   NOR2X1M U65 (.Y(\ab[6][4] ), 
	.B(n190), 
	.A(n35));
   NOR2X1M U66 (.Y(\ab[6][3] ), 
	.B(n190), 
	.A(n36));
   NOR2X1M U67 (.Y(\ab[6][2] ), 
	.B(n190), 
	.A(n37));
   NOR2X1M U68 (.Y(\ab[6][1] ), 
	.B(n190), 
	.A(n38));
   NOR2X1M U69 (.Y(\ab[6][0] ), 
	.B(n190), 
	.A(n39));
   NOR2X1M U70 (.Y(\ab[5][7] ), 
	.B(n191), 
	.A(n32));
   NOR2X1M U71 (.Y(\ab[5][6] ), 
	.B(n191), 
	.A(n173));
   NOR2X1M U72 (.Y(\ab[5][5] ), 
	.B(n191), 
	.A(n34));
   NOR2X1M U73 (.Y(\ab[5][4] ), 
	.B(n191), 
	.A(n35));
   NOR2X1M U74 (.Y(\ab[5][3] ), 
	.B(n191), 
	.A(n36));
   NOR2X1M U75 (.Y(\ab[5][2] ), 
	.B(n191), 
	.A(n37));
   NOR2X1M U76 (.Y(\ab[5][1] ), 
	.B(n191), 
	.A(n38));
   NOR2X1M U77 (.Y(\ab[5][0] ), 
	.B(n191), 
	.A(n39));
   NOR2X1M U78 (.Y(\ab[4][7] ), 
	.B(n192), 
	.A(n32));
   NOR2X1M U79 (.Y(\ab[4][6] ), 
	.B(n192), 
	.A(n173));
   NOR2X1M U80 (.Y(\ab[4][5] ), 
	.B(n192), 
	.A(n34));
   NOR2X1M U81 (.Y(\ab[4][4] ), 
	.B(n192), 
	.A(n35));
   NOR2X1M U82 (.Y(\ab[4][3] ), 
	.B(n192), 
	.A(n36));
   NOR2X1M U83 (.Y(\ab[4][2] ), 
	.B(n192), 
	.A(n37));
   NOR2X1M U84 (.Y(\ab[4][1] ), 
	.B(n192), 
	.A(n38));
   NOR2X1M U85 (.Y(\ab[4][0] ), 
	.B(n192), 
	.A(n39));
   NOR2X1M U86 (.Y(\ab[3][7] ), 
	.B(n193), 
	.A(n32));
   NOR2X1M U87 (.Y(\ab[3][6] ), 
	.B(n193), 
	.A(n173));
   NOR2X1M U88 (.Y(\ab[3][5] ), 
	.B(n193), 
	.A(n34));
   NOR2X1M U89 (.Y(\ab[3][4] ), 
	.B(n193), 
	.A(n35));
   NOR2X1M U90 (.Y(\ab[3][3] ), 
	.B(n193), 
	.A(n36));
   NOR2X1M U91 (.Y(\ab[3][2] ), 
	.B(n193), 
	.A(n37));
   NOR2X1M U92 (.Y(\ab[3][1] ), 
	.B(n193), 
	.A(n38));
   NOR2X1M U93 (.Y(\ab[3][0] ), 
	.B(n193), 
	.A(n39));
   NOR2X1M U94 (.Y(\ab[2][7] ), 
	.B(n194), 
	.A(n32));
   NOR2X1M U95 (.Y(\ab[2][6] ), 
	.B(n194), 
	.A(n173));
   NOR2X1M U96 (.Y(\ab[2][5] ), 
	.B(n194), 
	.A(n34));
   NOR2X1M U97 (.Y(\ab[2][4] ), 
	.B(n194), 
	.A(n35));
   NOR2X1M U98 (.Y(\ab[2][3] ), 
	.B(n194), 
	.A(n36));
   NOR2X1M U99 (.Y(\ab[2][2] ), 
	.B(n194), 
	.A(n37));
   NOR2X1M U100 (.Y(\ab[2][1] ), 
	.B(n194), 
	.A(n38));
   NOR2X1M U101 (.Y(\ab[2][0] ), 
	.B(n194), 
	.A(n39));
   NOR2X1M U102 (.Y(\ab[1][7] ), 
	.B(n30), 
	.A(n32));
   NOR2X1M U103 (.Y(\ab[1][6] ), 
	.B(n30), 
	.A(n173));
   NOR2X1M U104 (.Y(\ab[1][5] ), 
	.B(n30), 
	.A(n34));
   NOR2X1M U105 (.Y(\ab[1][4] ), 
	.B(n30), 
	.A(n35));
   NOR2X1M U106 (.Y(\ab[1][3] ), 
	.B(n30), 
	.A(n36));
   NOR2X1M U107 (.Y(\ab[1][2] ), 
	.B(n30), 
	.A(n37));
   NOR2X1M U108 (.Y(\ab[1][1] ), 
	.B(n30), 
	.A(n38));
   NOR2X1M U109 (.Y(\ab[1][0] ), 
	.B(n30), 
	.A(n39));
   NOR2X1M U110 (.Y(\ab[0][7] ), 
	.B(n31), 
	.A(n32));
   NOR2X1M U111 (.Y(\ab[0][6] ), 
	.B(n31), 
	.A(n173));
   NOR2X1M U112 (.Y(\ab[0][5] ), 
	.B(n31), 
	.A(n34));
   NOR2X1M U113 (.Y(\ab[0][4] ), 
	.B(n31), 
	.A(n35));
   NOR2X1M U114 (.Y(\ab[0][3] ), 
	.B(n31), 
	.A(n36));
   NOR2X1M U115 (.Y(\ab[0][2] ), 
	.B(n31), 
	.A(n37));
   NOR2X1M U116 (.Y(\ab[0][1] ), 
	.B(n31), 
	.A(n38));
   NOR2X1M U117 (.Y(PRODUCT[0]), 
	.B(n31), 
	.A(n39));
   ALU_00000008_00000004_DW01_add_1 FS_1 (.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }), 
	.B({ n10,
		n15,
		n16,
		n14,
		n13,
		n12,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }), 
	.CI(1'b0), 
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }));
endmodule

module ALU_00000008_00000004_test_1 (
	CLK, 
	RST_n, 
	A, 
	B, 
	ALU_FUN, 
	Enable, 
	ALU_OUT, 
	OUT_VALID, 
	test_si, 
	test_se, 
	FE_OFN12_RST_D1_M, 
	FE_OFN21_SE);
   input CLK;
   input RST_n;
   input [7:0] A;
   input [7:0] B;
   input [3:0] ALU_FUN;
   input Enable;
   output [15:0] ALU_OUT;
   output OUT_VALID;
   input test_si;
   input test_se;
   input FE_OFN12_RST_D1_M;
   input FE_OFN21_SE;

   // Internal wires
   wire N89;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N155;
   wire N156;
   wire N157;
   wire n10;
   wire n12;
   wire n15;
   wire n16;
   wire n17;
   wire n20;
   wire n21;
   wire n23;
   wire n24;
   wire n25;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n35;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n55;
   wire n56;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n128;
   wire n130;
   wire n132;
   wire n134;
   wire n136;
   wire n138;
   wire n140;
   wire n142;
   wire n144;
   wire n146;
   wire n148;
   wire n150;
   wire n152;
   wire n154;
   wire n156;
   wire n158;
   wire n160;
   wire n19;
   wire n22;
   wire n26;
   wire n27;
   wire n28;
   wire n34;
   wire n36;
   wire n42;
   wire n54;
   wire n57;
   wire n66;
   wire n75;
   wire n84;
   wire n93;
   wire n111;
   wire n117;
   wire n126;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;

   SDFFRQX2M \ALU_OUT_reg[8]  (.SI(ALU_OUT[7]), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(ALU_OUT[8]), 
	.D(n146), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[15]  (.SI(ALU_OUT[14]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(ALU_OUT[15]), 
	.D(n160), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[14]  (.SI(ALU_OUT[13]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(ALU_OUT[14]), 
	.D(n158), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[13]  (.SI(ALU_OUT[12]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(ALU_OUT[13]), 
	.D(n156), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[12]  (.SI(ALU_OUT[11]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(ALU_OUT[12]), 
	.D(n154), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[11]  (.SI(ALU_OUT[10]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(ALU_OUT[11]), 
	.D(n152), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[10]  (.SI(ALU_OUT[9]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(ALU_OUT[10]), 
	.D(n150), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[9]  (.SI(ALU_OUT[8]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(ALU_OUT[9]), 
	.D(n148), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[7]  (.SI(ALU_OUT[6]), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(ALU_OUT[7]), 
	.D(n144), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[6]  (.SI(ALU_OUT[5]), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(ALU_OUT[6]), 
	.D(n142), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[5]  (.SI(ALU_OUT[4]), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(ALU_OUT[5]), 
	.D(n140), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[4]  (.SI(ALU_OUT[3]), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(ALU_OUT[4]), 
	.D(n138), 
	.CK(CLK));
   SDFFRQX2M \ALU_OUT_reg[3]  (.SI(ALU_OUT[2]), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(ALU_OUT[3]), 
	.D(n136), 
	.CK(CLK));
   SDFFRHQX1M \ALU_OUT_reg[2]  (.SI(ALU_OUT[1]), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(ALU_OUT[2]), 
	.D(n134), 
	.CK(CLK));
   SDFFRHQX1M \ALU_OUT_reg[1]  (.SI(ALU_OUT[0]), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(ALU_OUT[1]), 
	.D(n132), 
	.CK(CLK));
   SDFFRHQX1M \ALU_OUT_reg[0]  (.SI(test_si), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(ALU_OUT[0]), 
	.D(n130), 
	.CK(CLK));
   SDFFRQX2M OUT_VALID_reg (.SI(ALU_OUT[15]), 
	.SE(FE_OFN21_SE), 
	.RN(RST_n), 
	.Q(OUT_VALID), 
	.D(n128), 
	.CK(CLK));
   NAND4X2M U3 (.Y(n24), 
	.D(n187), 
	.C(ALU_FUN[0]), 
	.B(Enable), 
	.A(n108));
   INVX2M U7 (.Y(n178), 
	.A(n103));
   NOR2BX2M U8 (.Y(n37), 
	.B(n187), 
	.AN(n102));
   NOR2X2M U9 (.Y(n12), 
	.B(n186), 
	.A(n185));
   NAND2X2M U10 (.Y(n44), 
	.B(n12), 
	.A(n32));
   NOR2BX2M U11 (.Y(n30), 
	.B(n33), 
	.AN(n32));
   NAND2X2M U12 (.Y(n103), 
	.B(n188), 
	.A(n38));
   NOR3X2M U13 (.Y(n32), 
	.C(n179), 
	.B(ALU_FUN[0]), 
	.A(n187));
   NOR3X2M U14 (.Y(n102), 
	.C(n179), 
	.B(ALU_FUN[3]), 
	.A(ALU_FUN[2]));
   NOR2X2M U15 (.Y(n108), 
	.B(ALU_FUN[3]), 
	.A(n186));
   NAND2X2M U16 (.Y(n33), 
	.B(n186), 
	.A(ALU_FUN[3]));
   INVX2M U17 (.Y(n177), 
	.A(n114));
   INVX2M U18 (.Y(n187), 
	.A(ALU_FUN[1]));
   INVX2M U19 (.Y(n181), 
	.A(n24));
   INVX2M U20 (.Y(n183), 
	.A(n106));
   INVX2M U21 (.Y(n188), 
	.A(ALU_FUN[0]));
   INVX2M U22 (.Y(n186), 
	.A(ALU_FUN[2]));
   INVX2M U23 (.Y(n185), 
	.A(ALU_FUN[3]));
   INVX2M U24 (.Y(n184), 
	.A(n107));
   NOR4X2M U26 (.Y(n25), 
	.D(ALU_FUN[1]), 
	.C(ALU_FUN[0]), 
	.B(n179), 
	.A(n33));
   NOR2BX2M U28 (.Y(n38), 
	.B(ALU_FUN[1]), 
	.AN(n102));
   INVX2M U29 (.Y(n180), 
	.A(n48));
   NOR2BX2M U30 (.Y(n115), 
	.B(ALU_FUN[3]), 
	.AN(n32));
   NOR2BX2M U31 (.Y(n29), 
	.B(ALU_FUN[0]), 
	.AN(n37));
   OAI22X1M U32 (.Y(n73), 
	.B1(n193), 
	.B0(n44), 
	.A1(n192), 
	.A0(n24));
   OAI22X1M U33 (.Y(n82), 
	.B1(n192), 
	.B0(n44), 
	.A1(n191), 
	.A0(n24));
   OAI22X1M U34 (.Y(n91), 
	.B1(n191), 
	.B0(n44), 
	.A1(n190), 
	.A0(n24));
   OAI22X1M U35 (.Y(n100), 
	.B1(n190), 
	.B0(n44), 
	.A1(n189), 
	.A0(n24));
   OAI22X1M U36 (.Y(n55), 
	.B1(n44), 
	.B0(n175), 
	.A1(n194), 
	.A0(n24));
   OAI22X1M U37 (.Y(n64), 
	.B1(n44), 
	.B0(n194), 
	.A1(n193), 
	.A0(n24));
   AOI222X4M U38 (.Y(n35), 
	.C1(n38), 
	.C0(N98), 
	.B1(n37), 
	.B0(N123), 
	.A1(n180), 
	.A0(A[1]));
   OAI222X2M U39 (.Y(n43), 
	.C1(n24), 
	.C0(n175), 
	.B1(n188), 
	.B0(n45), 
	.A1(n44), 
	.A0(n195));
   AOI221X2M U40 (.Y(n45), 
	.C0(n46), 
	.B1(n180), 
	.B0(A[2]), 
	.A1(n38), 
	.A0(N99));
   OAI2BB1X2M U41 (.Y(n46), 
	.B0(n47), 
	.A1N(n37), 
	.A0N(N124));
   NAND4BX1M U42 (.Y(n47), 
	.D(ALU_FUN[1]), 
	.C(Enable), 
	.B(N156), 
	.AN(n33));
   OAI21X2M U43 (.Y(n56), 
	.B0(n58), 
	.A1(n193), 
	.A0(n48));
   AOI22X1M U44 (.Y(n58), 
	.B1(n38), 
	.B0(N100), 
	.A1(n37), 
	.A0(N125));
   OAI21X2M U45 (.Y(n65), 
	.B0(n67), 
	.A1(n192), 
	.A0(n48));
   AOI22X1M U46 (.Y(n67), 
	.B1(n38), 
	.B0(N101), 
	.A1(n37), 
	.A0(N126));
   OAI21X2M U47 (.Y(n74), 
	.B0(n76), 
	.A1(n191), 
	.A0(n48));
   AOI22X1M U48 (.Y(n76), 
	.B1(n38), 
	.B0(N102), 
	.A1(n37), 
	.A0(N127));
   OAI21X2M U49 (.Y(n83), 
	.B0(n85), 
	.A1(n190), 
	.A0(n48));
   AOI22X1M U50 (.Y(n85), 
	.B1(n38), 
	.B0(N103), 
	.A1(n37), 
	.A0(N128));
   INVX2M U51 (.Y(n175), 
	.A(A[1]));
   AOI221XLM U52 (.Y(n60), 
	.C0(n183), 
	.B1(n194), 
	.B0(n184), 
	.A1(n25), 
	.A0(A[2]));
   AOI221XLM U53 (.Y(n69), 
	.C0(n183), 
	.B1(n193), 
	.B0(n184), 
	.A1(n25), 
	.A0(A[3]));
   AOI221XLM U54 (.Y(n78), 
	.C0(n183), 
	.B1(n192), 
	.B0(n184), 
	.A1(n25), 
	.A0(A[4]));
   AOI221XLM U55 (.Y(n87), 
	.C0(n183), 
	.B1(n191), 
	.B0(n184), 
	.A1(n25), 
	.A0(A[5]));
   AOI221XLM U56 (.Y(n96), 
	.C0(n183), 
	.B1(n190), 
	.B0(n184), 
	.A1(n25), 
	.A0(A[6]));
   AOI221XLM U57 (.Y(n105), 
	.C0(n183), 
	.B1(n189), 
	.B0(n184), 
	.A1(n25), 
	.A0(A[7]));
   AOI221XLM U58 (.Y(n50), 
	.C0(n183), 
	.B1(n175), 
	.B0(n184), 
	.A1(A[1]), 
	.A0(n25));
   AOI221XLM U59 (.Y(n49), 
	.C0(n181), 
	.B1(A[1]), 
	.B0(n182), 
	.A1(n175), 
	.A0(n25));
   AOI221XLM U60 (.Y(n59), 
	.C0(n181), 
	.B1(n182), 
	.B0(A[2]), 
	.A1(n194), 
	.A0(n25));
   AOI221XLM U61 (.Y(n68), 
	.C0(n181), 
	.B1(n182), 
	.B0(A[3]), 
	.A1(n193), 
	.A0(n25));
   AOI221XLM U62 (.Y(n77), 
	.C0(n181), 
	.B1(n182), 
	.B0(A[4]), 
	.A1(n192), 
	.A0(n25));
   AOI221XLM U63 (.Y(n86), 
	.C0(n181), 
	.B1(n182), 
	.B0(A[5]), 
	.A1(n191), 
	.A0(n25));
   AOI221XLM U64 (.Y(n95), 
	.C0(n181), 
	.B1(n182), 
	.B0(A[6]), 
	.A1(n190), 
	.A0(n25));
   AOI221XLM U65 (.Y(n104), 
	.C0(n181), 
	.B1(n182), 
	.B0(A[7]), 
	.A1(n189), 
	.A0(n25));
   NOR3BX2M U66 (.Y(n31), 
	.C(ALU_FUN[0]), 
	.B(n48), 
	.AN(N157));
   NAND3X2M U67 (.Y(n48), 
	.C(Enable), 
	.B(n187), 
	.A(n12));
   NAND4X2M U68 (.Y(n106), 
	.D(n188), 
	.C(ALU_FUN[1]), 
	.B(Enable), 
	.A(n108));
   NAND3X2M U69 (.Y(n107), 
	.C(n125), 
	.B(ALU_FUN[0]), 
	.A(Enable));
   AOI221XLM U70 (.Y(n125), 
	.C0(n12), 
	.B1(n185), 
	.B0(n187), 
	.A1(n186), 
	.A0(ALU_FUN[1]));
   INVX2M U71 (.Y(n179), 
	.A(Enable));
   OAI21X2M U72 (.Y(n92), 
	.B0(n94), 
	.A1(n189), 
	.A0(n48));
   AOI22X1M U73 (.Y(n94), 
	.B1(n38), 
	.B0(N104), 
	.A1(n37), 
	.A0(N129));
   NAND3X2M U74 (.Y(n114), 
	.C(n124), 
	.B(n106), 
	.A(n107));
   NAND3X2M U75 (.Y(n124), 
	.C(N106), 
	.B(ALU_FUN[0]), 
	.A(n38));
   INVX2M U76 (.Y(n182), 
	.A(n109));
   OAI211X2M U77 (.Y(n109), 
	.C0(Enable), 
	.B0(n187), 
	.A1(n110), 
	.A0(n108));
   NOR2X2M U78 (.Y(n110), 
	.B(n33), 
	.A(n188));
   AO22X1M U79 (.Y(n101), 
	.B1(n37), 
	.B0(N130), 
	.A1(n38), 
	.A0(N105));
   INVX2M U80 (.Y(n195), 
	.A(A[0]));
   INVX2M U81 (.Y(n190), 
	.A(A[6]));
   INVX2M U82 (.Y(n193), 
	.A(A[3]));
   INVX2M U83 (.Y(n192), 
	.A(A[4]));
   INVX2M U84 (.Y(n191), 
	.A(A[5]));
   INVX2M U85 (.Y(n189), 
	.A(A[7]));
   INVX2M U86 (.Y(n194), 
	.A(A[2]));
   NAND3X2M U88 (.Y(n130), 
	.C(n17), 
	.B(n16), 
	.A(n15));
   AOI221XLM U89 (.Y(n17), 
	.C0(n20), 
	.B1(n179), 
	.B0(ALU_OUT[0]), 
	.A1(n195), 
	.A0(n183));
   AOI221XLM U90 (.Y(n16), 
	.C0(n31), 
	.B1(N155), 
	.B0(n30), 
	.A1(n29), 
	.A0(N107));
   AOI2BB2X4M U91 (.Y(n15), 
	.B1(n178), 
	.B0(N89), 
	.A1N(n188), 
	.A0N(n35));
   NAND3BXLM U93 (.Y(n132), 
	.C(n41), 
	.B(n40), 
	.AN(n39));
   AOI221XLM U94 (.Y(n40), 
	.C0(n31), 
	.B1(n29), 
	.B0(N108), 
	.A1(n178), 
	.A0(N90));
   OAI2B2X1M U95 (.Y(n39), 
	.B1(n50), 
	.B0(B[1]), 
	.A1N(B[1]), 
	.A0(n49));
   AOI221X1M U96 (.Y(n41), 
	.C0(n43), 
	.B1(n179), 
	.B0(ALU_OUT[1]), 
	.A1(n175), 
	.A0(n183));
   NAND3BX2M U99 (.Y(n134), 
	.C(n53), 
	.B(n52), 
	.AN(n51));
   AOI221XLM U100 (.Y(n53), 
	.C0(n55), 
	.B1(n179), 
	.B0(ALU_OUT[2]), 
	.A1(n194), 
	.A0(n183));
   OAI2B2X1M U101 (.Y(n51), 
	.B1(n60), 
	.B0(B[2]), 
	.A1N(B[2]), 
	.A0(n59));
   AOI222X4M U102 (.Y(n52), 
	.C1(n178), 
	.C0(N91), 
	.B1(n29), 
	.B0(N109), 
	.A1(n56), 
	.A0(ALU_FUN[0]));
   NAND3BX2M U104 (.Y(n136), 
	.C(n63), 
	.B(n62), 
	.AN(n61));
   AOI221XLM U105 (.Y(n63), 
	.C0(n64), 
	.B1(n179), 
	.B0(ALU_OUT[3]), 
	.A1(n193), 
	.A0(n183));
   OAI2B2X1M U106 (.Y(n61), 
	.B1(n69), 
	.B0(B[3]), 
	.A1N(B[3]), 
	.A0(n68));
   AOI222X1M U107 (.Y(n62), 
	.C1(n178), 
	.C0(N92), 
	.B1(n29), 
	.B0(N110), 
	.A1(n65), 
	.A0(ALU_FUN[0]));
   NAND2X2M U109 (.Y(n160), 
	.B(n177), 
	.A(n123));
   AOI22X1M U110 (.Y(n123), 
	.B1(n179), 
	.B0(ALU_OUT[15]), 
	.A1(n115), 
	.A0(N122));
   NAND3BX2M U113 (.Y(n138), 
	.C(n72), 
	.B(n71), 
	.AN(n70));
   AOI221XLM U114 (.Y(n72), 
	.C0(n73), 
	.B1(n179), 
	.B0(ALU_OUT[4]), 
	.A1(n192), 
	.A0(n183));
   OAI2B2X1M U115 (.Y(n70), 
	.B1(n78), 
	.B0(B[4]), 
	.A1N(B[4]), 
	.A0(n77));
   AOI222X1M U116 (.Y(n71), 
	.C1(n178), 
	.C0(N93), 
	.B1(n29), 
	.B0(N111), 
	.A1(n74), 
	.A0(ALU_FUN[0]));
   NAND2X2M U117 (.Y(n158), 
	.B(n177), 
	.A(n122));
   AOI22X1M U118 (.Y(n122), 
	.B1(n179), 
	.B0(ALU_OUT[14]), 
	.A1(n115), 
	.A0(N121));
   NAND2X2M U119 (.Y(n154), 
	.B(n177), 
	.A(n120));
   AOI22X1M U120 (.Y(n120), 
	.B1(n179), 
	.B0(ALU_OUT[12]), 
	.A1(n115), 
	.A0(N119));
   NAND2X2M U121 (.Y(n156), 
	.B(n177), 
	.A(n121));
   AOI22X1M U122 (.Y(n121), 
	.B1(n179), 
	.B0(ALU_OUT[13]), 
	.A1(n115), 
	.A0(N120));
   NAND2X2M U123 (.Y(n150), 
	.B(n177), 
	.A(n118));
   AOI22X1M U124 (.Y(n118), 
	.B1(n179), 
	.B0(ALU_OUT[10]), 
	.A1(n115), 
	.A0(N117));
   NAND2X2M U125 (.Y(n152), 
	.B(n177), 
	.A(n119));
   AOI22X1M U126 (.Y(n119), 
	.B1(n179), 
	.B0(ALU_OUT[11]), 
	.A1(n115), 
	.A0(N118));
   INVX2M U127 (.Y(n173), 
	.A(B[6]));
   NAND3BX2M U128 (.Y(n144), 
	.C(n99), 
	.B(n98), 
	.AN(n97));
   AOI221XLM U129 (.Y(n99), 
	.C0(n100), 
	.B1(n179), 
	.B0(ALU_OUT[7]), 
	.A1(n189), 
	.A0(n183));
   OAI2B2X1M U130 (.Y(n97), 
	.B1(n105), 
	.B0(B[7]), 
	.A1N(B[7]), 
	.A0(n104));
   AOI222X1M U131 (.Y(n98), 
	.C1(n29), 
	.C0(N114), 
	.B1(n101), 
	.B0(ALU_FUN[0]), 
	.A1(n178), 
	.A0(N96));
   NAND2X2M U132 (.Y(n148), 
	.B(n177), 
	.A(n116));
   AOI22X1M U133 (.Y(n116), 
	.B1(n179), 
	.B0(ALU_OUT[9]), 
	.A1(n115), 
	.A0(N116));
   OAI2B11X2M U134 (.Y(n146), 
	.C0(n113), 
	.B0(n112), 
	.A1N(N97), 
	.A0(n103));
   AOI21X2M U135 (.Y(n113), 
	.B0(n114), 
	.A1(n179), 
	.A0(ALU_OUT[8]));
   AOI32X1M U136 (.Y(n112), 
	.B1(n115), 
	.B0(N115), 
	.A2(A[7]), 
	.A1(ALU_FUN[2]), 
	.A0(n32));
   INVX2M U137 (.Y(n176), 
	.A(n75));
   NAND3BX2M U138 (.Y(n140), 
	.C(n81), 
	.B(n80), 
	.AN(n79));
   AOI221XLM U139 (.Y(n81), 
	.C0(n82), 
	.B1(n179), 
	.B0(ALU_OUT[5]), 
	.A1(n191), 
	.A0(n183));
   OAI2B2X1M U157 (.Y(n79), 
	.B1(n87), 
	.B0(B[5]), 
	.A1N(B[5]), 
	.A0(n86));
   AOI222X1M U158 (.Y(n80), 
	.C1(n178), 
	.C0(N94), 
	.B1(n29), 
	.B0(N112), 
	.A1(n83), 
	.A0(ALU_FUN[0]));
   NAND3BX2M U159 (.Y(n142), 
	.C(n90), 
	.B(n89), 
	.AN(n88));
   AOI221XLM U160 (.Y(n90), 
	.C0(n91), 
	.B1(n179), 
	.B0(ALU_OUT[6]), 
	.A1(n190), 
	.A0(n183));
   OAI2B2X1M U161 (.Y(n88), 
	.B1(n96), 
	.B0(B[6]), 
	.A1N(B[6]), 
	.A0(n95));
   AOI222X1M U162 (.Y(n89), 
	.C1(n178), 
	.C0(N95), 
	.B1(n29), 
	.B0(N113), 
	.A1(n92), 
	.A0(ALU_FUN[0]));
   INVX2M U163 (.Y(n170), 
	.A(B[0]));
   OAI222X1M U164 (.Y(n20), 
	.C1(n24), 
	.C0(n195), 
	.B1(n23), 
	.B0(B[0]), 
	.A1(n170), 
	.A0(n21));
   AOI221XLM U165 (.Y(n21), 
	.C0(n181), 
	.B1(A[0]), 
	.B0(n182), 
	.A1(n195), 
	.A0(n25));
   AOI221XLM U166 (.Y(n23), 
	.C0(n183), 
	.B1(n195), 
	.B0(n184), 
	.A1(n25), 
	.A0(A[0]));
   INVX2M U167 (.Y(n174), 
	.A(n19));
   INVX2M U168 (.Y(n171), 
	.A(B[2]));
   INVX2M U169 (.Y(n172), 
	.A(B[3]));
   OAI2BB2X1M U170 (.Y(n128), 
	.B1(n179), 
	.B0(n10), 
	.A1N(n179), 
	.A0N(OUT_VALID));
   NOR3BX2M U171 (.Y(n10), 
	.C(n188), 
	.B(n187), 
	.AN(n12));
   NOR2X1M U172 (.Y(n166), 
	.B(B[7]), 
	.A(n189));
   NAND2BX1M U173 (.Y(n117), 
	.B(A[4]), 
	.AN(B[4]));
   NAND2BX1M U174 (.Y(n28), 
	.B(B[4]), 
	.AN(A[4]));
   CLKNAND2X2M U175 (.Y(n161), 
	.B(n28), 
	.A(n117));
   NOR2X1M U176 (.Y(n84), 
	.B(A[3]), 
	.A(n172));
   NOR2X1M U177 (.Y(n27), 
	.B(A[2]), 
	.A(n171));
   NOR2X1M U178 (.Y(n19), 
	.B(A[0]), 
	.A(n170));
   CLKNAND2X2M U179 (.Y(n111), 
	.B(n171), 
	.A(A[2]));
   NAND2BX1M U180 (.Y(n57), 
	.B(n111), 
	.AN(n27));
   AOI21X1M U181 (.Y(n22), 
	.B0(B[1]), 
	.A1(n175), 
	.A0(n19));
   AOI211X1M U182 (.Y(n26), 
	.C0(n22), 
	.B0(n57), 
	.A1(n174), 
	.A0(A[1]));
   CLKNAND2X2M U183 (.Y(n93), 
	.B(n172), 
	.A(A[3]));
   OAI31X1M U184 (.Y(n34), 
	.B0(n93), 
	.A2(n26), 
	.A1(n27), 
	.A0(n84));
   NAND2BX1M U185 (.Y(n164), 
	.B(B[5]), 
	.AN(A[5]));
   OAI211X1M U186 (.Y(n36), 
	.C0(n164), 
	.B0(n28), 
	.A1(n34), 
	.A0(n161));
   NAND2BX1M U187 (.Y(n126), 
	.B(A[5]), 
	.AN(B[5]));
   XNOR2X1M U188 (.Y(n163), 
	.B(B[6]), 
	.A(A[6]));
   AOI32X1M U189 (.Y(n42), 
	.B1(n190), 
	.B0(B[6]), 
	.A2(n163), 
	.A1(n126), 
	.A0(n36));
   CLKNAND2X2M U190 (.Y(n167), 
	.B(n189), 
	.A(B[7]));
   OAI21X1M U191 (.Y(N157), 
	.B0(n167), 
	.A1(n42), 
	.A0(n166));
   CLKNAND2X2M U192 (.Y(n66), 
	.B(n170), 
	.A(A[0]));
   OA21X1M U193 (.Y(n54), 
	.B0(B[1]), 
	.A1(n175), 
	.A0(n66));
   AOI211X1M U194 (.Y(n75), 
	.C0(n54), 
	.B0(n57), 
	.A1(n175), 
	.A0(n66));
   AOI31X1M U195 (.Y(n162), 
	.B0(n84), 
	.A2(n93), 
	.A1(n111), 
	.A0(n176));
   OAI2B11X1M U196 (.Y(n165), 
	.C0(n117), 
	.B0(n126), 
	.A1N(n162), 
	.A0(n161));
   AOI32X1M U197 (.Y(n168), 
	.B1(n173), 
	.B0(A[6]), 
	.A2(n163), 
	.A1(n164), 
	.A0(n165));
   AOI2B1X1M U198 (.Y(n169), 
	.B0(n166), 
	.A1N(n168), 
	.A0(n167));
   CLKINVX1M U199 (.Y(N156), 
	.A(n169));
   NOR2X1M U200 (.Y(N155), 
	.B(N156), 
	.A(N157));
   ALU_00000008_00000004_DW_div_uns_0 div_32 (.a({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.b({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.quotient({ N130,
		N129,
		N128,
		N127,
		N126,
		N125,
		N124,
		N123 }), 
	.n173(n173), 
	.n175(n175), 
	.n195(n195));
   ALU_00000008_00000004_DW01_sub_0 sub_30 (.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.CI(1'b0), 
	.DIFF({ N106,
		N105,
		N104,
		N103,
		N102,
		N101,
		N100,
		N99,
		N98 }), 
	.n170(n170), 
	.n173(n173), 
	.n172(n172), 
	.n195(n195), 
	.n171(n171));
   ALU_00000008_00000004_DW01_add_0 add_29 (.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.CI(1'b0), 
	.SUM({ N97,
		N96,
		N95,
		N94,
		N93,
		N92,
		N91,
		N90,
		N89 }));
   ALU_00000008_00000004_DW02_mult_0 mult_31 (.A({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }), 
	.B({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }), 
	.TC(1'b0), 
	.PRODUCT({ N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109,
		N108,
		N107 }), 
	.n170(n170), 
	.n172(n172), 
	.n189(n189), 
	.n190(n190), 
	.n175(n175), 
	.n195(n195), 
	.n171(n171), 
	.n191(n191), 
	.n192(n192), 
	.n193(n193), 
	.n194(n194), 
	.n173(n173));
endmodule

module UART_TX_test_1 (
	CLK, 
	RST_n, 
	P_DATA, 
	PAR_EN, 
	PAR_TYP, 
	DATA_VALID, 
	TX_OUT, 
	Busy, 
	test_si, 
	test_so, 
	test_se);
   input CLK;
   input RST_n;
   input [7:0] P_DATA;
   input PAR_EN;
   input PAR_TYP;
   input DATA_VALID;
   output TX_OUT;
   output Busy;
   input test_si;
   output test_so;
   input test_se;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire N25;
   wire N26;
   wire N27;
   wire N52;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n39;
   wire n40;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = n16 ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   SDFFRQX2M \Counter_reg[2]  (.SI(n39), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(N27), 
	.D(n37), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[0]  (.SI(N27), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[2]  (.SI(n15), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(current_state[2]), 
	.D(next_state[2]), 
	.CK(CLK));
   SDFFRQX2M \Counter_reg[1]  (.SI(n11), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(N26), 
	.D(n36), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[1]  (.SI(current_state[0]), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(current_state[1]), 
	.D(n9), 
	.CK(CLK));
   SDFFRQX2M \Counter_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(N25), 
	.D(n38), 
	.CK(CLK));
   INVX2M U9 (.Y(n10), 
	.A(n28));
   INVX2M U10 (.Y(n13), 
	.A(n27));
   NOR2X2M U11 (.Y(n28), 
	.B(Busy), 
	.A(DATA_VALID));
   AOI21X2M U12 (.Y(n24), 
	.B0(n28), 
	.A1(n13), 
	.A0(n11));
   OAI2B1X2M U13 (.Y(next_state[2]), 
	.B0(n10), 
	.A1N(n17), 
	.A0(n18));
   NAND2X2M U14 (.Y(n27), 
	.B(n23), 
	.A(n17));
   NAND2X2M U15 (.Y(Busy), 
	.B(n14), 
	.A(n20));
   INVX2M U16 (.Y(n12), 
	.A(n23));
   XOR3XLM U17 (.Y(n33), 
	.C(n34), 
	.B(P_DATA[0]), 
	.A(P_DATA[1]));
   XNOR2X2M U18 (.Y(n34), 
	.B(P_DATA[2]), 
	.A(P_DATA[3]));
   XOR3XLM U19 (.Y(n32), 
	.C(n35), 
	.B(P_DATA[4]), 
	.A(P_DATA[5]));
   XNOR2X2M U20 (.Y(n35), 
	.B(P_DATA[6]), 
	.A(P_DATA[7]));
   AOI211X2M U21 (.Y(n21), 
	.C0(current_state[1]), 
	.B0(current_state[0]), 
	.A1(n16), 
	.A0(n10));
   OAI31X1M U22 (.Y(next_state[0]), 
	.B0(n22), 
	.A2(n14), 
	.A1(n15), 
	.A0(n16));
   AOI31X2M U23 (.Y(n22), 
	.B0(n21), 
	.A2(n17), 
	.A1(n40), 
	.A0(n12));
   INVX2M U24 (.Y(n40), 
	.A(HTIE_LTIEHI_NET));
   OAI22X1M U25 (.Y(n36), 
	.B1(n25), 
	.B0(N26), 
	.A1(n39), 
	.A0(n24));
   OAI21X2M U26 (.Y(n37), 
	.B0(n26), 
	.A1(n25), 
	.A0(n39));
   OAI2BB1X2M U27 (.Y(n26), 
	.B0(N27), 
	.A1N(n24), 
	.A0N(n27));
   INVX2M U28 (.Y(n9), 
	.A(n19));
   AOI221XLM U29 (.Y(n19), 
	.C0(n21), 
	.B1(current_state[0]), 
	.B0(n20), 
	.A1(n17), 
	.A0(n18));
   OAI22X1M U30 (.Y(n38), 
	.B1(n27), 
	.B0(N25), 
	.A1(n10), 
	.A0(n11));
   NOR3X2M U31 (.Y(n17), 
	.C(n15), 
	.B(current_state[2]), 
	.A(current_state[0]));
   NOR2X2M U32 (.Y(n20), 
	.B(current_state[1]), 
	.A(current_state[2]));
   NAND3X2M U33 (.Y(n23), 
	.C(N27), 
	.B(N25), 
	.A(N26));
   NAND2X2M U34 (.Y(n25), 
	.B(N25), 
	.A(n13));
   INVX2M U35 (.Y(n11), 
	.A(N25));
   INVX2M U36 (.Y(n15), 
	.A(current_state[1]));
   INVX2M U37 (.Y(n14), 
	.A(current_state[0]));
   INVX2M U38 (.Y(n39), 
	.A(N26));
   INVX2M U39 (.Y(n16), 
	.A(current_state[2]));
   NAND2X2M U40 (.Y(n18), 
	.B(n12), 
	.A(HTIE_LTIEHI_NET));
   OAI211X2M U41 (.Y(TX_OUT), 
	.C0(n30), 
	.B0(Busy), 
	.A1(n16), 
	.A0(n29));
   NOR2X2M U42 (.Y(n29), 
	.B(n31), 
	.A(current_state[1]));
   AOI2BB2XLM U43 (.Y(n30), 
	.B1(current_state[1]), 
	.B0(N52), 
	.A1N(n20), 
	.A0N(n14));
   XOR3XLM U44 (.Y(n31), 
	.C(n33), 
	.B(n32), 
	.A(LTIE_LTIELO_NET));
   MX2X2M U45 (.Y(N52), 
	.S0(N27), 
	.B(n7), 
	.A(n8));
   MX4X1M U46 (.Y(n7), 
	.S1(N26), 
	.S0(N25), 
	.D(P_DATA[7]), 
	.C(P_DATA[6]), 
	.B(P_DATA[5]), 
	.A(P_DATA[4]));
   MX4X1M U47 (.Y(n8), 
	.S1(N26), 
	.S0(N25), 
	.D(P_DATA[3]), 
	.C(P_DATA[2]), 
	.B(P_DATA[1]), 
	.A(P_DATA[0]));
endmodule

module data_sampling_10_test_1 (
	CLK, 
	RST_n, 
	RX_IN, 
	Prescale, 
	data_samp_en, 
	edge_cnt, 
	sampled_bit, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN22_SE);
   input CLK;
   input RST_n;
   input RX_IN;
   input [5:0] Prescale;
   input data_samp_en;
   input [3:0] edge_cnt;
   output sampled_bit;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN22_SE;

   // Internal wires
   wire first_value;
   wire second_value;
   wire third_value;
   wire out_next_1;
   wire out_next_2;
   wire out_next_3;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n8;

   assign test_so = out_next_3 ;

   SDFFRQX2M out_next_2_reg (.SI(out_next_1), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(out_next_2), 
	.D(second_value), 
	.CK(CLK));
   SDFFRQX2M out_next_1_reg (.SI(test_si), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(out_next_1), 
	.D(first_value), 
	.CK(CLK));
   SDFFRQX2M out_next_3_reg (.SI(out_next_2), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(out_next_3), 
	.D(third_value), 
	.CK(CLK));
   OAI2B2X1M U6 (.Y(sampled_bit), 
	.B1(n16), 
	.B0(n3), 
	.A1N(first_value), 
	.A0(n15));
   INVX2M U7 (.Y(n1), 
	.A(n19));
   NOR4BX1M U8 (.Y(n19), 
	.D(n18), 
	.C(edge_cnt[2]), 
	.B(edge_cnt[1]), 
	.AN(n20));
   NOR2X2M U9 (.Y(n20), 
	.B(n4), 
	.A(n2));
   INVX2M U10 (.Y(n2), 
	.A(data_samp_en));
   NOR4X1M U11 (.Y(n18), 
	.D(edge_cnt[2]), 
	.C(edge_cnt[1]), 
	.B(edge_cnt[0]), 
	.A(n4));
   INVX2M U12 (.Y(n4), 
	.A(edge_cnt[3]));
   INVX2M U13 (.Y(n3), 
	.A(second_value));
   NOR2BX2M U14 (.Y(n16), 
	.B(first_value), 
	.AN(n15));
   AOI22X1M U15 (.Y(n15), 
	.B1(n19), 
	.B0(RX_IN), 
	.A1(out_next_3), 
	.A0(n1));
   OAI2BB2X1M U16 (.Y(first_value), 
	.B1(n21), 
	.B0(n8), 
	.A1N(n21), 
	.A0N(out_next_1));
   NAND4X2M U17 (.Y(n21), 
	.D(edge_cnt[0]), 
	.C(n22), 
	.B(edge_cnt[1]), 
	.A(edge_cnt[2]));
   NOR2X2M U18 (.Y(n22), 
	.B(n2), 
	.A(edge_cnt[3]));
   OAI2BB2X1M U19 (.Y(second_value), 
	.B1(n17), 
	.B0(n8), 
	.A1N(n17), 
	.A0N(out_next_2));
   NAND2X2M U20 (.Y(n17), 
	.B(data_samp_en), 
	.A(n18));
   OAI2BB2X1M U21 (.Y(third_value), 
	.B1(n8), 
	.B0(n13), 
	.A1N(out_next_3), 
	.A0N(n13));
   NAND4X2M U22 (.Y(n13), 
	.D(data_samp_en), 
	.C(n14), 
	.B(edge_cnt[0]), 
	.A(edge_cnt[3]));
   NOR2X2M U23 (.Y(n14), 
	.B(edge_cnt[1]), 
	.A(edge_cnt[2]));
   INVX2M U24 (.Y(n8), 
	.A(RX_IN));
endmodule

module edge_bit_counter_10_test_1 (
	CLK, 
	RST_n, 
	parity_en, 
	enable, 
	bit_cnt, 
	edge_cnt, 
	test_si, 
	test_so, 
	test_se);
   input CLK;
   input RST_n;
   input parity_en;
   input enable;
   output [3:0] bit_cnt;
   output [3:0] edge_cnt;
   input test_si;
   output test_so;
   input test_se;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire \add_37/carry[4] ;
   wire \add_37/carry[3] ;
   wire \add_37/carry[2] ;
   wire n14;
   wire n15;
   wire n16;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n46;
   wire [3:0] Bit_Counter;
   wire [4:0] Edge_Counter;

   assign test_so = n24 ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRQX2M \Edge_Counter_reg[4]  (.SI(Edge_Counter[3]), 
	.SE(test_se), 
	.RN(n14), 
	.Q(Edge_Counter[4]), 
	.D(n43), 
	.CK(CLK));
   SDFFRQX2M \Bit_Counter_reg[3]  (.SI(n25), 
	.SE(test_se), 
	.RN(n14), 
	.Q(Bit_Counter[3]), 
	.D(n44), 
	.CK(CLK));
   SDFFRQX2M \Bit_Counter_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(n14), 
	.Q(Bit_Counter[0]), 
	.D(n45), 
	.CK(CLK));
   SDFFRQX2M \Bit_Counter_reg[2]  (.SI(Bit_Counter[1]), 
	.SE(test_se), 
	.RN(n14), 
	.Q(Bit_Counter[2]), 
	.D(n41), 
	.CK(CLK));
   SDFFRQX2M \Bit_Counter_reg[1]  (.SI(n22), 
	.SE(test_se), 
	.RN(n14), 
	.Q(Bit_Counter[1]), 
	.D(n42), 
	.CK(CLK));
   SDFFRX1M \Edge_Counter_reg[0]  (.SI(n23), 
	.SE(test_se), 
	.RN(RST_n), 
	.QN(n20), 
	.Q(Edge_Counter[0]), 
	.D(n40), 
	.CK(CLK));
   SDFFRX1M \Edge_Counter_reg[3]  (.SI(Edge_Counter[2]), 
	.SE(test_se), 
	.RN(n14), 
	.QN(n17), 
	.Q(Edge_Counter[3]), 
	.D(n37), 
	.CK(CLK));
   SDFFRX1M \Edge_Counter_reg[2]  (.SI(Edge_Counter[1]), 
	.SE(test_se), 
	.RN(n14), 
	.QN(n18), 
	.Q(Edge_Counter[2]), 
	.D(n38), 
	.CK(CLK));
   SDFFRX1M \Edge_Counter_reg[1]  (.SI(Edge_Counter[0]), 
	.SE(test_se), 
	.RN(n14), 
	.QN(n19), 
	.Q(Edge_Counter[1]), 
	.D(n39), 
	.CK(CLK));
   NOR2X2M U16 (.Y(bit_cnt[0]), 
	.B(n22), 
	.A(n15));
   INVX2M U17 (.Y(n21), 
	.A(n28));
   INVX2M U18 (.Y(n16), 
	.A(n32));
   INVX2M U19 (.Y(n14), 
	.A(n15));
   INVX2M U20 (.Y(n15), 
	.A(RST_n));
   NOR2X2M U21 (.Y(bit_cnt[1]), 
	.B(n46), 
	.A(n15));
   NOR2X2M U22 (.Y(bit_cnt[2]), 
	.B(n25), 
	.A(n15));
   NOR2X2M U23 (.Y(bit_cnt[3]), 
	.B(n23), 
	.A(n15));
   NAND2X2M U24 (.Y(n28), 
	.B(n33), 
	.A(enable));
   NAND2X2M U25 (.Y(n32), 
	.B(n24), 
	.A(enable));
   NOR2X2M U26 (.Y(edge_cnt[1]), 
	.B(n19), 
	.A(n15));
   NOR2X2M U27 (.Y(edge_cnt[2]), 
	.B(n18), 
	.A(n15));
   NOR2X2M U28 (.Y(edge_cnt[0]), 
	.B(n20), 
	.A(n15));
   NOR2X2M U29 (.Y(edge_cnt[3]), 
	.B(n17), 
	.A(n15));
   INVX2M U30 (.Y(n46), 
	.A(Bit_Counter[1]));
   INVX2M U31 (.Y(n25), 
	.A(Bit_Counter[2]));
   NAND3BX2M U32 (.Y(n26), 
	.C(enable), 
	.B(Edge_Counter[4]), 
	.AN(n33));
   OAI32X1M U33 (.Y(n42), 
	.B1(n46), 
	.B0(n31), 
	.A2(n22), 
	.A1(Bit_Counter[1]), 
	.A0(n28));
   AOI21X2M U34 (.Y(n31), 
	.B0(n16), 
	.A1(n22), 
	.A0(n21));
   OAI32X1M U35 (.Y(n41), 
	.B1(n25), 
	.B0(n30), 
	.A2(n29), 
	.A1(Bit_Counter[2]), 
	.A0(n28));
   AOI21X2M U36 (.Y(n30), 
	.B0(n16), 
	.A1(n29), 
	.A0(n21));
   OAI22X1M U37 (.Y(n44), 
	.B1(n28), 
	.B0(n34), 
	.A1(n32), 
	.A0(n23));
   AOI2BB1X2M U38 (.Y(n34), 
	.B0(Bit_Counter[3]), 
	.A1N(n25), 
	.A0N(n29));
   OAI22X1M U39 (.Y(n45), 
	.B1(n28), 
	.B0(Bit_Counter[0]), 
	.A1(n32), 
	.A0(n22));
   NOR2BX2M U40 (.Y(n27), 
	.B(Edge_Counter[4]), 
	.AN(enable));
   OAI2BB2X1M U41 (.Y(n37), 
	.B1(n17), 
	.B0(n26), 
	.A1N(n27), 
	.A0N(N18));
   OAI2BB2X1M U42 (.Y(n38), 
	.B1(n18), 
	.B0(n26), 
	.A1N(n27), 
	.A0N(N17));
   OAI2BB2X1M U43 (.Y(n39), 
	.B1(n19), 
	.B0(n26), 
	.A1N(n27), 
	.A0N(N16));
   OAI2B2X1M U44 (.Y(n40), 
	.B1(n20), 
	.B0(n26), 
	.A1N(n27), 
	.A0(Edge_Counter[0]));
   OAI2BB1X2M U45 (.Y(n43), 
	.B0(n26), 
	.A1N(n27), 
	.A0N(N19));
   INVX2M U46 (.Y(n22), 
	.A(Bit_Counter[0]));
   INVX2M U47 (.Y(n23), 
	.A(Bit_Counter[3]));
   OAI32X1M U48 (.Y(n33), 
	.B1(n24), 
	.B0(n36), 
	.A2(Bit_Counter[1]), 
	.A1(Bit_Counter[2]), 
	.A0(n35));
   AOI31X2M U49 (.Y(n36), 
	.B0(n23), 
	.A2(n22), 
	.A1(n25), 
	.A0(n46));
   NAND2X2M U50 (.Y(n35), 
	.B(Edge_Counter[4]), 
	.A(HTIE_LTIEHI_NET));
   NAND2X2M U51 (.Y(n29), 
	.B(Bit_Counter[0]), 
	.A(Bit_Counter[1]));
   INVX2M U52 (.Y(n24), 
	.A(Edge_Counter[4]));
   ADDHX1M U53 (.S(N16), 
	.CO(\add_37/carry[2] ), 
	.B(Edge_Counter[0]), 
	.A(Edge_Counter[1]));
   ADDHX1M U54 (.S(N17), 
	.CO(\add_37/carry[3] ), 
	.B(\add_37/carry[2] ), 
	.A(Edge_Counter[2]));
   ADDHX1M U55 (.S(N18), 
	.CO(\add_37/carry[4] ), 
	.B(\add_37/carry[3] ), 
	.A(Edge_Counter[3]));
   CLKXOR2X2M U56 (.Y(N19), 
	.B(Edge_Counter[4]), 
	.A(\add_37/carry[4] ));
endmodule

module Parity_Check (
	par_typ, 
	par_chk_en, 
	sampled_bit, 
	p_data, 
	par_err);
   input par_typ;
   input par_chk_en;
   input sampled_bit;
   input [7:0] p_data;
   output par_err;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;

   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   XOR3XLM U2 (.Y(n1), 
	.C(n4), 
	.B(n3), 
	.A(n2));
   XOR3XLM U3 (.Y(n3), 
	.C(n5), 
	.B(p_data[4]), 
	.A(p_data[5]));
   XOR3XLM U4 (.Y(n2), 
	.C(n6), 
	.B(p_data[0]), 
	.A(p_data[1]));
   XNOR2X2M U5 (.Y(n4), 
	.B(LTIE_LTIELO_NET), 
	.A(sampled_bit));
   NOR2BX2M U6 (.Y(par_err), 
	.B(n1), 
	.AN(par_chk_en));
   XNOR2X2M U7 (.Y(n6), 
	.B(p_data[2]), 
	.A(p_data[3]));
   XNOR2X2M U8 (.Y(n5), 
	.B(p_data[6]), 
	.A(p_data[7]));
endmodule

module Start_Check_test_1 (
	CLK, 
	RST_n, 
	strt_chk_en, 
	sampled_bit, 
	strt_glitch, 
	test_si, 
	test_se);
   input CLK;
   input RST_n;
   input strt_chk_en;
   input sampled_bit;
   output strt_glitch;
   input test_si;
   input test_se;

   // Internal wires
   wire n2;

   SDFFRQX2M strt_glitch_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(strt_glitch), 
	.D(n2), 
	.CK(CLK));
   AO2B2X2M U2 (.Y(n2), 
	.B1(sampled_bit), 
	.B0(strt_chk_en), 
	.A1N(strt_chk_en), 
	.A0(strt_glitch));
endmodule

module Stop_Check_test_1 (
	CLK, 
	RST_n, 
	stp_chk_en, 
	sampled_bit, 
	stp_err, 
	test_si, 
	test_se);
   input CLK;
   input RST_n;
   input stp_chk_en;
   input sampled_bit;
   output stp_err;
   input test_si;
   input test_se;

   // Internal wires
   wire N5;

   SDFFRQX2M stp_err_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(stp_err), 
	.D(N5), 
	.CK(CLK));
   NOR2BX2M U4 (.Y(N5), 
	.B(sampled_bit), 
	.AN(stp_chk_en));
endmodule

module deserializer_test_1 (
	CLK, 
	RST_n, 
	deser_en, 
	bit_cnt, 
	sampled_bit, 
	P_DATA, 
	test_si, 
	test_se, 
	FE_OFN14_RST_D2_M, 
	FE_OFN18_SE, 
	FE_OFN22_SE);
   input CLK;
   input RST_n;
   input deser_en;
   input [3:0] bit_cnt;
   input sampled_bit;
   output [7:0] P_DATA;
   input test_si;
   input test_se;
   input FE_OFN14_RST_D2_M;
   input FE_OFN18_SE;
   input FE_OFN22_SE;

   // Internal wires
   wire \index[0] ;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n1;
   wire n2;
   wire n11;

   assign \index[0]  = bit_cnt[0] ;

   SDFFRQX2M \P_DATA_reg[5]  (.SI(P_DATA[4]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(P_DATA[5]), 
	.D(n35), 
	.CK(CLK));
   SDFFRQX2M \P_DATA_reg[1]  (.SI(P_DATA[0]), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN14_RST_D2_M), 
	.Q(P_DATA[1]), 
	.D(n31), 
	.CK(CLK));
   SDFFRQX2M \P_DATA_reg[4]  (.SI(P_DATA[3]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(P_DATA[4]), 
	.D(n34), 
	.CK(CLK));
   SDFFRQX2M \P_DATA_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(FE_OFN14_RST_D2_M), 
	.Q(P_DATA[0]), 
	.D(n30), 
	.CK(CLK));
   SDFFRQX2M \P_DATA_reg[7]  (.SI(P_DATA[6]), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(P_DATA[7]), 
	.D(n37), 
	.CK(CLK));
   SDFFRQX2M \P_DATA_reg[3]  (.SI(P_DATA[2]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(P_DATA[3]), 
	.D(n33), 
	.CK(CLK));
   SDFFRQX2M \P_DATA_reg[6]  (.SI(P_DATA[5]), 
	.SE(FE_OFN22_SE), 
	.RN(RST_n), 
	.Q(P_DATA[6]), 
	.D(n36), 
	.CK(CLK));
   SDFFRQX2M \P_DATA_reg[2]  (.SI(P_DATA[1]), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(P_DATA[2]), 
	.D(n32), 
	.CK(CLK));
   INVX2M U11 (.Y(n11), 
	.A(n20));
   INVX2M U12 (.Y(n2), 
	.A(n15));
   NOR2BX2M U13 (.Y(n16), 
	.B(\index[0] ), 
	.AN(n25));
   NOR2X2M U14 (.Y(n27), 
	.B(bit_cnt[1]), 
	.A(\index[0] ));
   CLKXOR2X2M U15 (.Y(n20), 
	.B(\index[0] ), 
	.A(bit_cnt[1]));
   AND2X2M U16 (.Y(n18), 
	.B(n25), 
	.A(\index[0] ));
   CLKXOR2X2M U17 (.Y(n15), 
	.B(bit_cnt[2]), 
	.A(n27));
   INVX2M U18 (.Y(n1), 
	.A(sampled_bit));
   AND2X2M U19 (.Y(n25), 
	.B(deser_en), 
	.A(n28));
   CLKXOR2X2M U20 (.Y(n28), 
	.B(bit_cnt[3]), 
	.A(n29));
   NAND2BX2M U21 (.Y(n29), 
	.B(n27), 
	.AN(bit_cnt[2]));
   OAI2BB2X1M U22 (.Y(n30), 
	.B1(n1), 
	.B0(n14), 
	.A1N(n14), 
	.A0N(P_DATA[0]));
   NAND3X2M U23 (.Y(n14), 
	.C(n16), 
	.B(n15), 
	.A(n11));
   OAI2BB2X1M U24 (.Y(n31), 
	.B1(n17), 
	.B0(n1), 
	.A1N(n17), 
	.A0N(P_DATA[1]));
   NAND3X2M U25 (.Y(n17), 
	.C(n18), 
	.B(n15), 
	.A(n11));
   OAI2BB2X1M U26 (.Y(n32), 
	.B1(n19), 
	.B0(n1), 
	.A1N(n19), 
	.A0N(P_DATA[2]));
   NAND3X2M U27 (.Y(n19), 
	.C(n16), 
	.B(n20), 
	.A(n15));
   OAI2BB2X1M U28 (.Y(n33), 
	.B1(n21), 
	.B0(n1), 
	.A1N(n21), 
	.A0N(P_DATA[3]));
   NAND3X2M U29 (.Y(n21), 
	.C(n18), 
	.B(n20), 
	.A(n15));
   OAI2BB2X1M U30 (.Y(n34), 
	.B1(n22), 
	.B0(n1), 
	.A1N(n22), 
	.A0N(P_DATA[4]));
   NAND3X2M U31 (.Y(n22), 
	.C(n2), 
	.B(n16), 
	.A(n11));
   OAI2BB2X1M U32 (.Y(n35), 
	.B1(n23), 
	.B0(n1), 
	.A1N(n23), 
	.A0N(P_DATA[5]));
   NAND3X2M U33 (.Y(n23), 
	.C(n2), 
	.B(n18), 
	.A(n11));
   OAI2BB2X1M U34 (.Y(n36), 
	.B1(n24), 
	.B0(n1), 
	.A1N(n24), 
	.A0N(P_DATA[6]));
   NAND3X2M U35 (.Y(n24), 
	.C(n2), 
	.B(n20), 
	.A(n16));
   OAI2BB2X1M U36 (.Y(n37), 
	.B1(n26), 
	.B0(n1), 
	.A1N(n26), 
	.A0N(P_DATA[7]));
   NAND3X2M U37 (.Y(n26), 
	.C(n2), 
	.B(n20), 
	.A(n18));
endmodule

module UART_RX_10_test_1 (
	CLK, 
	RST_n, 
	PAR_TYP, 
	PAR_EN, 
	Prescale, 
	RX_IN, 
	P_DATA, 
	DATA_Valid, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN14_RST_D2_M, 
	FE_OFN18_SE, 
	FE_OFN22_SE);
   input CLK;
   input RST_n;
   input PAR_TYP;
   input PAR_EN;
   input [5:0] Prescale;
   input RX_IN;
   output [7:0] P_DATA;
   output DATA_Valid;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN14_RST_D2_M;
   input FE_OFN18_SE;
   input FE_OFN22_SE;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire sampled_bit;
   wire enable;
   wire par_chk_en;
   wire par_err;
   wire strt_chk_en;
   wire strt_glitch;
   wire stp_err;
   wire deser_en;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N75;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N179;
   wire N180;
   wire N181;
   wire N182;
   wire N183;
   wire N184;
   wire N185;
   wire N186;
   wire n43;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire \r113/EQ ;
   wire \add_202/carry[3] ;
   wire \r112/carry[2] ;
   wire \r112/carry[3] ;
   wire n1;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n41;
   wire n42;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire [3:0] edge_cnt;
   wire [3:0] bit_cnt;
   wire [7:0] p_data;
   wire [3:0] middle_sample_point;
   wire [2:0] current_state;
   wire [2:0] next_state;
   wire [7:0] out_next;

   assign test_so = stp_err ;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   SDFFRQX2M \out_next_reg[7]  (.SI(out_next[6]), 
	.SE(test_se), 
	.RN(FE_OFN14_RST_D2_M), 
	.Q(out_next[7]), 
	.D(P_DATA[7]), 
	.CK(CLK));
   SDFFRQX2M \out_next_reg[6]  (.SI(out_next[5]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(out_next[6]), 
	.D(P_DATA[6]), 
	.CK(CLK));
   SDFFRQX2M \out_next_reg[5]  (.SI(out_next[4]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(out_next[5]), 
	.D(P_DATA[5]), 
	.CK(CLK));
   SDFFRQX2M \out_next_reg[4]  (.SI(out_next[3]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(out_next[4]), 
	.D(P_DATA[4]), 
	.CK(CLK));
   SDFFRQX2M \out_next_reg[3]  (.SI(out_next[2]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(out_next[3]), 
	.D(P_DATA[3]), 
	.CK(CLK));
   SDFFRQX2M \out_next_reg[2]  (.SI(out_next[1]), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(out_next[2]), 
	.D(P_DATA[2]), 
	.CK(CLK));
   SDFFRQX2M \out_next_reg[1]  (.SI(out_next[0]), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(out_next[1]), 
	.D(P_DATA[1]), 
	.CK(CLK));
   SDFFRQX2M \out_next_reg[0]  (.SI(n88), 
	.SE(test_se), 
	.RN(FE_OFN14_RST_D2_M), 
	.Q(out_next[0]), 
	.D(P_DATA[0]), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[2]  (.SI(n85), 
	.SE(test_se), 
	.RN(FE_OFN14_RST_D2_M), 
	.Q(current_state[2]), 
	.D(next_state[2]), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(FE_OFN14_RST_D2_M), 
	.Q(current_state[0]), 
	.D(next_state[0]), 
	.CK(CLK));
   SDFFRQX2M \current_state_reg[1]  (.SI(n83), 
	.SE(test_se), 
	.RN(FE_OFN14_RST_D2_M), 
	.Q(current_state[1]), 
	.D(next_state[1]), 
	.CK(CLK));
   NOR2X2M U4 (.Y(n1), 
	.B(n9), 
	.A(current_state[1]));
   OAI211X2M U8 (.Y(enable), 
	.C0(n82), 
	.B0(n62), 
	.A1(n76), 
	.A0(n83));
   INVX2M U9 (.Y(n51), 
	.A(n67));
   NAND2X2M U10 (.Y(n61), 
	.B(n53), 
	.A(n84));
   INVX2M U11 (.Y(n53), 
	.A(N102));
   NOR3BX2M U12 (.Y(n59), 
	.C(bit_cnt[2]), 
	.B(bit_cnt[1]), 
	.AN(\r113/EQ ));
   INVX2M U21 (.Y(n84), 
	.A(n78));
   NAND3BX2M U22 (.Y(n68), 
	.C(n59), 
	.B(n81), 
	.AN(bit_cnt[3]));
   NAND3X2M U23 (.Y(n67), 
	.C(bit_cnt[3]), 
	.B(n81), 
	.A(n59));
   NOR3BX2M U24 (.Y(n58), 
	.C(n62), 
	.B(bit_cnt[2]), 
	.AN(bit_cnt[3]));
   NAND3X2M U25 (.Y(n64), 
	.C(n73), 
	.B(bit_cnt[3]), 
	.A(bit_cnt[0]));
   NOR3X2M U26 (.Y(n73), 
	.C(bit_cnt[1]), 
	.B(bit_cnt[2]), 
	.A(N75));
   INVX2M U27 (.Y(n81), 
	.A(bit_cnt[0]));
   NAND2X2M U28 (.Y(n66), 
	.B(n64), 
	.A(n60));
   INVX2M U29 (.Y(N79), 
	.A(middle_sample_point[1]));
   INVX2M U30 (.Y(n52), 
	.A(n79));
   NOR3X2M U31 (.Y(DATA_Valid), 
	.C(n78), 
	.B(n83), 
	.A(n79));
   NAND2X2M U32 (.Y(n78), 
	.B(n85), 
	.A(current_state[2]));
   NAND2X2M U33 (.Y(n62), 
	.B(n83), 
	.A(n84));
   INVX2M U34 (.Y(n43), 
	.A(n55));
   OAI211X2M U35 (.Y(n55), 
	.C0(\r113/EQ ), 
	.B0(n58), 
	.A1(n57), 
	.A0(n56));
   NOR3X2M U36 (.Y(n60), 
	.C(n85), 
	.B(current_state[2]), 
	.A(n83));
   NAND3X2M U37 (.Y(next_state[2]), 
	.C(n63), 
	.B(n62), 
	.A(n61));
   AOI32X1M U38 (.Y(n63), 
	.B1(n60), 
	.B0(n50), 
	.A2(deser_en), 
	.A1(n86), 
	.A0(n51));
   INVX2M U39 (.Y(n50), 
	.A(n64));
   NOR3BX2M U40 (.Y(n56), 
	.C(bit_cnt[0]), 
	.B(n86), 
	.AN(bit_cnt[1]));
   OAI21X2M U41 (.Y(middle_sample_point[1]), 
	.B0(n75), 
	.A1(n87), 
	.A0(N78));
   NAND2X2M U43 (.Y(n75), 
	.B(N78), 
	.A(n87));
   INVX2M U44 (.Y(n82), 
	.A(n77));
   NAND2X2M U45 (.Y(n76), 
	.B(n85), 
	.A(n53));
   AOI31X2M U46 (.Y(n77), 
	.B0(current_state[2]), 
	.A2(n83), 
	.A1(n85), 
	.A0(RX_IN));
   MX2X2M U47 (.Y(P_DATA[0]), 
	.S0(n1), 
	.B(n10), 
	.A(out_next[0]));
   AND2X2M U48 (.Y(n10), 
	.B(current_state[2]), 
	.A(N179));
   AO22X1M U49 (.Y(N179), 
	.B1(n52), 
	.B0(p_data[0]), 
	.A1(n79), 
	.A0(out_next[0]));
   MX2X2M U50 (.Y(P_DATA[1]), 
	.S0(n1), 
	.B(n11), 
	.A(out_next[1]));
   AND2X2M U51 (.Y(n11), 
	.B(current_state[2]), 
	.A(N180));
   AO22X1M U52 (.Y(N180), 
	.B1(n52), 
	.B0(p_data[1]), 
	.A1(n79), 
	.A0(out_next[1]));
   MX2X2M U53 (.Y(P_DATA[2]), 
	.S0(n1), 
	.B(n12), 
	.A(out_next[2]));
   AND2X2M U54 (.Y(n12), 
	.B(current_state[2]), 
	.A(N181));
   AO22X1M U55 (.Y(N181), 
	.B1(n52), 
	.B0(p_data[2]), 
	.A1(n79), 
	.A0(out_next[2]));
   MX2X2M U56 (.Y(P_DATA[3]), 
	.S0(n1), 
	.B(n13), 
	.A(out_next[3]));
   AND2X2M U57 (.Y(n13), 
	.B(current_state[2]), 
	.A(N182));
   AO22X1M U58 (.Y(N182), 
	.B1(n52), 
	.B0(p_data[3]), 
	.A1(n79), 
	.A0(out_next[3]));
   MX2X2M U59 (.Y(P_DATA[4]), 
	.S0(n1), 
	.B(n14), 
	.A(out_next[4]));
   AND2X2M U60 (.Y(n14), 
	.B(current_state[2]), 
	.A(N183));
   AO22X1M U61 (.Y(N183), 
	.B1(n52), 
	.B0(p_data[4]), 
	.A1(n79), 
	.A0(out_next[4]));
   MX2X2M U62 (.Y(P_DATA[5]), 
	.S0(n1), 
	.B(n15), 
	.A(out_next[5]));
   AND2X2M U63 (.Y(n15), 
	.B(current_state[2]), 
	.A(N184));
   AO22X1M U64 (.Y(N184), 
	.B1(n52), 
	.B0(p_data[5]), 
	.A1(n79), 
	.A0(out_next[5]));
   MX2X2M U65 (.Y(P_DATA[6]), 
	.S0(n1), 
	.B(n16), 
	.A(out_next[6]));
   AND2X2M U66 (.Y(n16), 
	.B(current_state[2]), 
	.A(N185));
   AO22X1M U67 (.Y(N185), 
	.B1(n52), 
	.B0(p_data[6]), 
	.A1(n79), 
	.A0(out_next[6]));
   MX2X2M U68 (.Y(P_DATA[7]), 
	.S0(n1), 
	.B(n17), 
	.A(out_next[7]));
   AND2X2M U69 (.Y(n17), 
	.B(current_state[2]), 
	.A(N186));
   AO22X1M U70 (.Y(N186), 
	.B1(n52), 
	.B0(p_data[7]), 
	.A1(n79), 
	.A0(out_next[7]));
   NAND2X2M U71 (.Y(n79), 
	.B(n80), 
	.A(N102));
   OAI33X2M U72 (.Y(n80), 
	.B2(stp_err), 
	.B1(strt_glitch), 
	.B0(par_err), 
	.A2(stp_err), 
	.A1(strt_glitch), 
	.A0(HTIE_LTIEHI_NET));
   AND4X2M U73 (.Y(par_chk_en), 
	.D(n60), 
	.C(bit_cnt[0]), 
	.B(bit_cnt[3]), 
	.A(n59));
   INVX2M U74 (.Y(n83), 
	.A(current_state[0]));
   INVX2M U76 (.Y(n85), 
	.A(current_state[1]));
   OAI31X1M U77 (.Y(n71), 
	.B0(n66), 
	.A2(current_state[1]), 
	.A1(current_state[2]), 
	.A0(n72));
   AOI2BB2XLM U78 (.Y(n72), 
	.B1(n68), 
	.B0(current_state[0]), 
	.A1N(current_state[0]), 
	.A0N(RX_IN));
   OAI221X1M U79 (.Y(next_state[0]), 
	.C0(n70), 
	.B1(n61), 
	.B0(n83), 
	.A1(n54), 
	.A0(n69));
   INVX2M U80 (.Y(n54), 
	.A(n58));
   AOI22X1M U81 (.Y(n69), 
	.B1(\r113/EQ ), 
	.B0(n56), 
	.A1(n57), 
	.A0(N83));
   AOI31X2M U82 (.Y(n70), 
	.B0(n71), 
	.A2(deser_en), 
	.A1(HTIE_LTIEHI_NET), 
	.A0(n51));
   NOR4X1M U83 (.Y(strt_chk_en), 
	.D(current_state[2]), 
	.C(current_state[1]), 
	.B(n68), 
	.A(n83));
   OAI2B11X2M U84 (.Y(next_state[1]), 
	.C0(n66), 
	.B0(n65), 
	.A1N(strt_chk_en), 
	.A0(strt_glitch));
   OAI21X2M U85 (.Y(n65), 
	.B0(deser_en), 
	.A1(n67), 
	.A0(HTIE_LTIEHI_NET));
   NOR3X2M U86 (.Y(deser_en), 
	.C(n85), 
	.B(current_state[2]), 
	.A(current_state[0]));
   XNOR2X2M U87 (.Y(n9), 
	.B(n18), 
	.A(current_state[0]));
   INVX2M U88 (.Y(n18), 
	.A(current_state[2]));
   NOR3X2M U89 (.Y(n57), 
	.C(n81), 
	.B(bit_cnt[1]), 
	.A(HTIE_LTIEHI_NET));
   XNOR2X2M U90 (.Y(middle_sample_point[2]), 
	.B(n75), 
	.A(LTIE_LTIELO_NET));
   CLKXOR2X2M U91 (.Y(middle_sample_point[3]), 
	.B(n74), 
	.A(HTIE_LTIEHI_NET));
   NOR2X2M U92 (.Y(n74), 
	.B(n75), 
	.A(LTIE_LTIELO_NET));
   INVX2M U93 (.Y(n87), 
	.A(LTIE_LTIELO_NET));
   INVX2M U94 (.Y(n86), 
	.A(HTIE_LTIEHI_NET));
   INVX2M U95 (.Y(N78), 
	.A(LTIE_LTIELO_NET));
   OR2X2M U96 (.Y(n5), 
	.B(LTIE_LTIELO_NET), 
	.A(LTIE_LTIELO_NET));
   AND2X1M U97 (.Y(N82), 
	.B(middle_sample_point[3]), 
	.A(\add_202/carry[3] ));
   CLKXOR2X2M U98 (.Y(N81), 
	.B(\add_202/carry[3] ), 
	.A(middle_sample_point[3]));
   AND2X1M U99 (.Y(\add_202/carry[3] ), 
	.B(middle_sample_point[2]), 
	.A(middle_sample_point[1]));
   CLKXOR2X2M U100 (.Y(N80), 
	.B(middle_sample_point[1]), 
	.A(middle_sample_point[2]));
   AND2X1M U101 (.Y(N50), 
	.B(middle_sample_point[3]), 
	.A(\r112/carry[3] ));
   CLKXOR2X2M U102 (.Y(N49), 
	.B(\r112/carry[3] ), 
	.A(middle_sample_point[3]));
   AND2X1M U103 (.Y(\r112/carry[3] ), 
	.B(middle_sample_point[2]), 
	.A(\r112/carry[2] ));
   CLKXOR2X2M U104 (.Y(N48), 
	.B(\r112/carry[2] ), 
	.A(middle_sample_point[2]));
   OR2X1M U105 (.Y(\r112/carry[2] ), 
	.B(N78), 
	.A(middle_sample_point[1]));
   XNOR2X1M U106 (.Y(N47), 
	.B(middle_sample_point[1]), 
	.A(N78));
   CLKINVX1M U107 (.Y(N95), 
	.A(LTIE_LTIELO_NET));
   OAI2BB1X1M U108 (.Y(N96), 
	.B0(n5), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(LTIE_LTIELO_NET));
   OR2X1M U109 (.Y(n6), 
	.B(LTIE_LTIELO_NET), 
	.A(n5));
   OAI2BB1X1M U110 (.Y(N97), 
	.B0(n6), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(n5));
   OR2X1M U111 (.Y(n7), 
	.B(LTIE_LTIELO_NET), 
	.A(n6));
   OAI2BB1X1M U112 (.Y(N98), 
	.B0(n7), 
	.A1N(LTIE_LTIELO_NET), 
	.A0N(n6));
   OR2X1M U113 (.Y(n8), 
	.B(HTIE_LTIEHI_NET), 
	.A(n7));
   OAI2BB1X1M U114 (.Y(N99), 
	.B0(n8), 
	.A1N(HTIE_LTIEHI_NET), 
	.A0N(n7));
   NOR2X1M U115 (.Y(N101), 
	.B(LTIE_LTIELO_NET), 
	.A(n8));
   AO21XLM U116 (.Y(N100), 
	.B0(N101), 
	.A1(LTIE_LTIELO_NET), 
	.A0(n8));
   NOR2BX1M U117 (.Y(n19), 
	.B(edge_cnt[0]), 
	.AN(LTIE_LTIELO_NET));
   OAI2B2X1M U118 (.Y(n25), 
	.B1(n19), 
	.B0(N47), 
	.A1N(edge_cnt[1]), 
	.A0(n19));
   NOR2BX1M U119 (.Y(n20), 
	.B(LTIE_LTIELO_NET), 
	.AN(edge_cnt[0]));
   OAI2B2X1M U120 (.Y(n24), 
	.B1(n20), 
	.B0(edge_cnt[1]), 
	.A1N(N47), 
	.A0(n20));
   CLKXOR2X2M U121 (.Y(n22), 
	.B(edge_cnt[3]), 
	.A(N49));
   CLKXOR2X2M U122 (.Y(n21), 
	.B(edge_cnt[2]), 
	.A(N48));
   NOR2X1M U123 (.Y(n23), 
	.B(n21), 
	.A(n22));
   NAND4BX1M U124 (.Y(N75), 
	.D(n23), 
	.C(n24), 
	.B(n25), 
	.AN(N50));
   CLKINVX1M U125 (.Y(\r113/EQ ), 
	.A(N75));
   XNOR2X1M U126 (.Y(n44), 
	.B(edge_cnt[2]), 
	.A(N97));
   NOR2BX1M U127 (.Y(n26), 
	.B(edge_cnt[0]), 
	.AN(N95));
   OAI2B2X1M U128 (.Y(n42), 
	.B1(n26), 
	.B0(N96), 
	.A1N(edge_cnt[1]), 
	.A0(n26));
   XNOR2X1M U129 (.Y(n41), 
	.B(edge_cnt[3]), 
	.A(N98));
   NOR2BX1M U130 (.Y(n27), 
	.B(N95), 
	.AN(edge_cnt[0]));
   OAI2B2X1M U131 (.Y(n28), 
	.B1(n27), 
	.B0(edge_cnt[1]), 
	.A1N(N96), 
	.A0(n27));
   NOR4BX1M U132 (.Y(n29), 
	.D(N99), 
	.C(N100), 
	.B(N101), 
	.AN(n28));
   AND4X1M U133 (.Y(N102), 
	.D(n29), 
	.C(n41), 
	.B(n42), 
	.A(n44));
   XNOR2X1M U134 (.Y(n46), 
	.B(edge_cnt[2]), 
	.A(N80));
   XNOR2X1M U135 (.Y(n45), 
	.B(edge_cnt[3]), 
	.A(N81));
   CLKNAND2X2M U136 (.Y(n49), 
	.B(n45), 
	.A(n46));
   CLKXOR2X2M U137 (.Y(n48), 
	.B(edge_cnt[1]), 
	.A(N79));
   CLKXOR2X2M U138 (.Y(n47), 
	.B(edge_cnt[0]), 
	.A(N78));
   NOR4X1M U139 (.Y(N83), 
	.D(n47), 
	.C(N82), 
	.B(n48), 
	.A(n49));
   data_sampling_10_test_1 dut_sample (.CLK(CLK), 
	.RST_n(RST_n), 
	.RX_IN(RX_IN), 
	.Prescale({ Prescale[5],
		Prescale[4],
		Prescale[3],
		Prescale[2],
		Prescale[1],
		Prescale[0] }), 
	.data_samp_en(enable), 
	.edge_cnt({ edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }), 
	.sampled_bit(sampled_bit), 
	.test_si(p_data[7]), 
	.test_so(n89), 
	.test_se(test_se), 
	.FE_OFN22_SE(FE_OFN22_SE));
   edge_bit_counter_10_test_1 edge_bit_dut (.CLK(CLK), 
	.RST_n(RST_n), 
	.parity_en(PAR_EN), 
	.enable(enable), 
	.bit_cnt({ bit_cnt[3],
		bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }), 
	.edge_cnt({ edge_cnt[3],
		edge_cnt[2],
		edge_cnt[1],
		edge_cnt[0] }), 
	.test_si(n89), 
	.test_so(n88), 
	.test_se(test_se));
   Parity_Check parity_dut (.par_typ(PAR_TYP), 
	.par_chk_en(par_chk_en), 
	.sampled_bit(sampled_bit), 
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }), 
	.par_err(par_err));
   Start_Check_test_1 srt_dut (.CLK(CLK), 
	.RST_n(FE_OFN14_RST_D2_M), 
	.strt_chk_en(strt_chk_en), 
	.sampled_bit(sampled_bit), 
	.strt_glitch(strt_glitch), 
	.test_si(out_next[7]), 
	.test_se(test_se));
   Stop_Check_test_1 stp_dut (.CLK(CLK), 
	.RST_n(FE_OFN14_RST_D2_M), 
	.stp_chk_en(n43), 
	.sampled_bit(sampled_bit), 
	.stp_err(stp_err), 
	.test_si(strt_glitch), 
	.test_se(test_se));
   deserializer_test_1 deser_dut (.CLK(CLK), 
	.RST_n(RST_n), 
	.deser_en(deser_en), 
	.bit_cnt({ bit_cnt[3],
		bit_cnt[2],
		bit_cnt[1],
		bit_cnt[0] }), 
	.sampled_bit(sampled_bit), 
	.P_DATA({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }), 
	.test_si(n18), 
	.test_se(test_se), 
	.FE_OFN14_RST_D2_M(FE_OFN14_RST_D2_M), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.FE_OFN22_SE(FE_OFN22_SE));
endmodule

module Bit_Sync_00000002_00000005_test_1 (
	RST_n, 
	CLK, 
	ASYNC, 
	SYNC, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN18_SE);
   input RST_n;
   input CLK;
   input [4:0] ASYNC;
   output [4:0] SYNC;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN18_SE;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire \FF_Stage[1][4] ;
   wire \FF_Stage[1][3] ;
   wire \FF_Stage[1][2] ;
   wire \FF_Stage[1][1] ;
   wire \FF_Stage[1][0] ;
   wire \FF_Stage[0][4] ;
   wire \FF_Stage[0][3] ;
   wire \FF_Stage[0][2] ;
   wire \FF_Stage[0][1] ;
   wire \FF_Stage[0][0] ;

   assign test_so2 = \FF_Stage[1][4]  ;
   assign test_so1 = \FF_Stage[0][2]  ;

   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   SDFFRQX2M \FF_Stage_reg[1][4]  (.SI(\FF_Stage[1][3] ), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][4] ), 
	.D(\FF_Stage[0][4] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][3]  (.SI(\FF_Stage[1][2] ), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][3] ), 
	.D(\FF_Stage[0][3] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][2]  (.SI(\FF_Stage[1][1] ), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][2] ), 
	.D(\FF_Stage[0][2] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][1]  (.SI(\FF_Stage[1][0] ), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][1] ), 
	.D(\FF_Stage[0][1] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][0]  (.SI(\FF_Stage[0][4] ), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][0] ), 
	.D(\FF_Stage[0][0] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][4]  (.SI(\FF_Stage[0][3] ), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][4] ), 
	.D(LTIE_LTIELO_NET), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][3]  (.SI(test_si2), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][3] ), 
	.D(ASYNC[3]), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][2]  (.SI(\FF_Stage[0][1] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][2] ), 
	.D(ASYNC[2]), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][1]  (.SI(\FF_Stage[0][0] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][1] ), 
	.D(ASYNC[1]), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][0]  (.SI(test_si1), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][0] ), 
	.D(ASYNC[0]), 
	.CK(CLK));
   AND2X2M U13 (.Y(SYNC[0]), 
	.B(RST_n), 
	.A(\FF_Stage[1][0] ));
   AND2X2M U14 (.Y(SYNC[1]), 
	.B(RST_n), 
	.A(\FF_Stage[1][1] ));
   AND2X2M U15 (.Y(SYNC[4]), 
	.B(RST_n), 
	.A(\FF_Stage[1][4] ));
   AND2X2M U16 (.Y(SYNC[3]), 
	.B(RST_n), 
	.A(\FF_Stage[1][3] ));
   AND2X2M U17 (.Y(SYNC[2]), 
	.B(RST_n), 
	.A(\FF_Stage[1][2] ));
endmodule

module Bit_Sync_00000002_00000005_test_0 (
	RST_n, 
	CLK, 
	ASYNC, 
	SYNC, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN17_SE, 
	FE_OFN18_SE);
   input RST_n;
   input CLK;
   input [4:0] ASYNC;
   output [4:0] SYNC;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN17_SE;
   input FE_OFN18_SE;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire \FF_Stage[1][4] ;
   wire \FF_Stage[1][3] ;
   wire \FF_Stage[1][2] ;
   wire \FF_Stage[1][1] ;
   wire \FF_Stage[1][0] ;
   wire \FF_Stage[0][4] ;
   wire \FF_Stage[0][3] ;
   wire \FF_Stage[0][2] ;
   wire \FF_Stage[0][1] ;
   wire \FF_Stage[0][0] ;

   assign test_so = \FF_Stage[1][4]  ;

   TIELOM LTIE_LTIELO (.Y(LTIE_LTIELO_NET));
   SDFFRQX2M \FF_Stage_reg[1][4]  (.SI(\FF_Stage[1][3] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][4] ), 
	.D(\FF_Stage[0][4] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][0]  (.SI(\FF_Stage[0][4] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][0] ), 
	.D(\FF_Stage[0][0] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][3]  (.SI(\FF_Stage[1][2] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][3] ), 
	.D(\FF_Stage[0][3] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][2]  (.SI(\FF_Stage[1][1] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][2] ), 
	.D(\FF_Stage[0][2] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[1][1]  (.SI(\FF_Stage[1][0] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[1][1] ), 
	.D(\FF_Stage[0][1] ), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][4]  (.SI(\FF_Stage[0][3] ), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][4] ), 
	.D(LTIE_LTIELO_NET), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][3]  (.SI(\FF_Stage[0][2] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][3] ), 
	.D(ASYNC[3]), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][2]  (.SI(\FF_Stage[0][1] ), 
	.SE(FE_OFN17_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][2] ), 
	.D(ASYNC[2]), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][1]  (.SI(\FF_Stage[0][0] ), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][1] ), 
	.D(ASYNC[1]), 
	.CK(CLK));
   SDFFRQX2M \FF_Stage_reg[0][0]  (.SI(test_si), 
	.SE(FE_OFN18_SE), 
	.RN(RST_n), 
	.Q(\FF_Stage[0][0] ), 
	.D(ASYNC[0]), 
	.CK(CLK));
   AND2X2M U13 (.Y(SYNC[0]), 
	.B(RST_n), 
	.A(\FF_Stage[1][0] ));
   AND2X2M U14 (.Y(SYNC[3]), 
	.B(RST_n), 
	.A(\FF_Stage[1][3] ));
   AND2X2M U15 (.Y(SYNC[1]), 
	.B(RST_n), 
	.A(\FF_Stage[1][1] ));
   AND2X2M U16 (.Y(SYNC[2]), 
	.B(RST_n), 
	.A(\FF_Stage[1][2] ));
   AND2X2M U17 (.Y(SYNC[4]), 
	.B(RST_n), 
	.A(\FF_Stage[1][4] ));
endmodule

module fifo_wrptr_full_00000008_00000010_test_1 (
	W_CLK, 
	W_RST, 
	W_INC, 
	gray_Rptr, 
	WFULL, 
	Waddr, 
	gray_Wptr, 
	test_si, 
	test_se, 
	FE_OFN11_RST_D1_M, 
	FE_OFN12_RST_D1_M, 
	FE_OFN18_SE, 
	FE_OFN21_SE, 
	REF_CLK_M__L5_N2);
   input W_CLK;
   input W_RST;
   input W_INC;
   input [4:0] gray_Rptr;
   output WFULL;
   output [3:0] Waddr;
   output [4:0] gray_Wptr;
   input test_si;
   input test_se;
   input FE_OFN11_RST_D1_M;
   input FE_OFN12_RST_D1_M;
   input FE_OFN18_SE;
   input FE_OFN21_SE;
   input REF_CLK_M__L5_N2;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N116;
   wire n4;
   wire n6;
   wire n8;
   wire n10;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n22;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n31;
   wire n33;
   wire n35;
   wire n37;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire \add_59/carry[4] ;
   wire \add_59/carry[3] ;
   wire \add_59/carry[2] ;
   wire n9;
   wire n11;
   wire n21;
   wire n23;
   wire n29;
   wire n50;
   wire n51;
   wire [4:0] Wptr;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRQX2M \gray_Wptr_reg[3]  (.SI(gray_Wptr[2]), 
	.SE(FE_OFN18_SE), 
	.RN(W_RST), 
	.Q(gray_Wptr[3]), 
	.D(n37), 
	.CK(W_CLK));
   SDFFRQX2M \gray_Wptr_reg[2]  (.SI(gray_Wptr[1]), 
	.SE(FE_OFN18_SE), 
	.RN(W_RST), 
	.Q(gray_Wptr[2]), 
	.D(n35), 
	.CK(W_CLK));
   SDFFRQX2M \gray_Wptr_reg[1]  (.SI(gray_Wptr[0]), 
	.SE(FE_OFN18_SE), 
	.RN(W_RST), 
	.Q(gray_Wptr[1]), 
	.D(n33), 
	.CK(W_CLK));
   SDFFRQX2M \gray_Wptr_reg[0]  (.SI(n43), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(gray_Wptr[0]), 
	.D(n31), 
	.CK(W_CLK));
   SDFFRQX2M \Wptr_reg[3]  (.SI(n50), 
	.SE(test_se), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(N116), 
	.D(n45), 
	.CK(W_CLK));
   SDFFRQX2M \Wptr_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(Wptr[0]), 
	.D(n49), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \Wptr_reg[2]  (.SI(Wptr[1]), 
	.SE(test_se), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(Wptr[2]), 
	.D(n46), 
	.CK(W_CLK));
   SDFFRX1M \Wptr_reg[4]  (.SI(n51), 
	.SE(FE_OFN18_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.QN(n43), 
	.Q(Wptr[4]), 
	.D(n48), 
	.CK(W_CLK));
   SDFFRX1M \Wptr_reg[1]  (.SI(Wptr[0]), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.QN(n44), 
	.Q(Wptr[1]), 
	.D(n47), 
	.CK(REF_CLK_M__L5_N2));
   NOR2X3M U7 (.Y(Waddr[2]), 
	.B(n9), 
	.A(n50));
   INVX2M U8 (.Y(n21), 
	.A(n26));
   CLKINVX2M U9 (.Y(n9), 
	.A(FE_OFN12_RST_D1_M));
   AOI22X1M U10 (.Y(n26), 
	.B1(n20), 
	.B0(n23), 
	.A1(gray_Rptr[1]), 
	.A0(n28));
   XNOR2X2M U11 (.Y(n28), 
	.B(gray_Rptr[3]), 
	.A(gray_Rptr[2]));
   CLKXOR2X2M U12 (.Y(n20), 
	.B(gray_Rptr[3]), 
	.A(gray_Rptr[2]));
   INVX2M U13 (.Y(n23), 
	.A(gray_Rptr[1]));
   NOR2X4M U14 (.Y(Waddr[3]), 
	.B(n9), 
	.A(n51));
   OAI2BB2X1M U15 (.Y(n45), 
	.B1(n51), 
	.B0(n10), 
	.A1N(n10), 
	.A0N(N44));
   OAI2BB2X1M U16 (.Y(n46), 
	.B1(n50), 
	.B0(n10), 
	.A1N(n10), 
	.A0N(N43));
   INVX2M U17 (.Y(n11), 
	.A(gray_Rptr[4]));
   NOR2BX2M U19 (.Y(n10), 
	.B(WFULL), 
	.AN(W_INC));
   NOR2X2M U20 (.Y(Waddr[0]), 
	.B(n9), 
	.A(n29));
   OAI2B2X1M U21 (.Y(n16), 
	.B1(n26), 
	.B0(gray_Rptr[0]), 
	.A1N(gray_Rptr[0]), 
	.A0(n27));
   AOI22X1M U22 (.Y(n27), 
	.B1(n23), 
	.B0(n28), 
	.A1(n20), 
	.A0(gray_Rptr[1]));
   AOI22X1M U23 (.Y(n24), 
	.B1(n16), 
	.B0(n44), 
	.A1(n21), 
	.A0(n25));
   NAND2BX2M U24 (.Y(n25), 
	.B(Wptr[0]), 
	.AN(n16));
   AND4X2M U25 (.Y(WFULL), 
	.D(n14), 
	.C(n13), 
	.B(Wptr[4]), 
	.A(n12));
   NAND3X2M U26 (.Y(n13), 
	.C(n44), 
	.B(n11), 
	.A(n21));
   AOI211X2M U27 (.Y(n14), 
	.C0(n18), 
	.B0(n17), 
	.A1(n16), 
	.A0(n15));
   OAI2BB2X1M U28 (.Y(n12), 
	.B1(n24), 
	.B0(gray_Rptr[4]), 
	.A1N(n44), 
	.A0N(n29));
   XNOR2X2M U29 (.Y(n18), 
	.B(n19), 
	.A(Wptr[2]));
   NAND2X2M U30 (.Y(n19), 
	.B(n11), 
	.A(n20));
   XNOR2X2M U31 (.Y(n17), 
	.B(n22), 
	.A(N116));
   NAND2X2M U32 (.Y(n22), 
	.B(n11), 
	.A(gray_Rptr[3]));
   OAI2BB2X1M U33 (.Y(n47), 
	.B1(n10), 
	.B0(n44), 
	.A1N(n10), 
	.A0N(N42));
   OAI2B2X1M U34 (.Y(n49), 
	.B1(n29), 
	.B0(n10), 
	.A1N(n10), 
	.A0(Wptr[0]));
   OAI2BB2X1M U35 (.Y(n48), 
	.B1(n10), 
	.B0(n43), 
	.A1N(n10), 
	.A0N(N45));
   INVX2M U36 (.Y(n29), 
	.A(Wptr[0]));
   INVX2M U37 (.Y(n50), 
	.A(Wptr[2]));
   INVX2M U38 (.Y(n51), 
	.A(N116));
   NOR2X2M U39 (.Y(n15), 
	.B(Wptr[0]), 
	.A(gray_Rptr[4]));
   NOR2X2M U40 (.Y(Waddr[1]), 
	.B(n9), 
	.A(n44));
   OAI2BB2X1M U41 (.Y(n33), 
	.B1(n6), 
	.B0(Wptr[4]), 
	.A1N(Wptr[4]), 
	.A0N(gray_Wptr[1]));
   XNOR2X2M U42 (.Y(n6), 
	.B(n50), 
	.A(n44));
   OAI2BB2X1M U43 (.Y(n35), 
	.B1(Wptr[4]), 
	.B0(n8), 
	.A1N(Wptr[4]), 
	.A0N(gray_Wptr[2]));
   XNOR2X2M U54 (.Y(n8), 
	.B(Wptr[2]), 
	.A(N116));
   OAI2BB2X1M U55 (.Y(n37), 
	.B1(n51), 
	.B0(Wptr[4]), 
	.A1N(Wptr[4]), 
	.A0N(gray_Wptr[3]));
   OAI2BB2X1M U56 (.Y(n31), 
	.B1(n4), 
	.B0(Wptr[4]), 
	.A1N(Wptr[4]), 
	.A0N(gray_Wptr[0]));
   XNOR2X2M U57 (.Y(n4), 
	.B(n29), 
	.A(n44));
   ADDHX1M U58 (.S(N43), 
	.CO(\add_59/carry[3] ), 
	.B(\add_59/carry[2] ), 
	.A(Wptr[2]));
   ADDHX1M U59 (.S(N42), 
	.CO(\add_59/carry[2] ), 
	.B(Wptr[0]), 
	.A(Wptr[1]));
   ADDHX1M U60 (.S(N44), 
	.CO(\add_59/carry[4] ), 
	.B(\add_59/carry[3] ), 
	.A(N116));
   CLKXOR2X2M U61 (.Y(N45), 
	.B(Wptr[4]), 
	.A(\add_59/carry[4] ));
   INVX2M U3 (.Y(gray_Wptr[4]), 
	.A(HTIE_LTIEHI_NET));
endmodule

module fifo_rdptr_empty_00000008_00000010_test_1 (
	R_CLK, 
	R_RST, 
	R_INC, 
	gray_Wptr, 
	REMPTY, 
	Raddr, 
	gray_Rptr, 
	test_si, 
	test_se, 
	FE_OFN18_SE, 
	FE_OFN24_SE);
   input R_CLK;
   input R_RST;
   input R_INC;
   input [4:0] gray_Wptr;
   output REMPTY;
   output [3:0] Raddr;
   output [4:0] gray_Rptr;
   input test_si;
   input test_se;
   input FE_OFN18_SE;
   input FE_OFN24_SE;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire N41;
   wire N42;
   wire N43;
   wire N44;
   wire N115;
   wire n3;
   wire n4;
   wire n5;
   wire n7;
   wire n11;
   wire n13;
   wire n17;
   wire n19;
   wire n21;
   wire n23;
   wire n25;
   wire n27;
   wire n29;
   wire n31;
   wire n33;
   wire \eq_41/A[1] ;
   wire \add_65/carry[4] ;
   wire \add_65/carry[3] ;
   wire \add_65/carry[2] ;
   wire n6;
   wire n8;
   wire n9;
   wire n10;
   wire n12;
   wire n14;
   wire n15;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire [4:0] Rptr;
   wire [3:0] Wptr;

   TIEHIM HTIE_LTIEHI (.Y(HTIE_LTIEHI_NET));
   SDFFRQX2M \gray_Rptr_reg[3]  (.SI(gray_Rptr[2]), 
	.SE(FE_OFN18_SE), 
	.RN(R_RST), 
	.Q(gray_Rptr[3]), 
	.D(n23), 
	.CK(R_CLK));
   SDFFRQX2M \gray_Rptr_reg[2]  (.SI(gray_Rptr[1]), 
	.SE(FE_OFN18_SE), 
	.RN(R_RST), 
	.Q(gray_Rptr[2]), 
	.D(n21), 
	.CK(R_CLK));
   SDFFRQX2M \gray_Rptr_reg[1]  (.SI(gray_Rptr[0]), 
	.SE(test_se), 
	.RN(R_RST), 
	.Q(gray_Rptr[1]), 
	.D(n19), 
	.CK(R_CLK));
   SDFFRQX2M \gray_Rptr_reg[0]  (.SI(Rptr[4]), 
	.SE(test_se), 
	.RN(R_RST), 
	.Q(gray_Rptr[0]), 
	.D(n17), 
	.CK(R_CLK));
   SDFFRQX2M \Rptr_reg[0]  (.SI(test_si), 
	.SE(test_se), 
	.RN(R_RST), 
	.Q(Rptr[0]), 
	.D(n33), 
	.CK(R_CLK));
   SDFFRQX2M \Rptr_reg[3]  (.SI(n37), 
	.SE(FE_OFN24_SE), 
	.RN(R_RST), 
	.Q(N115), 
	.D(n25), 
	.CK(R_CLK));
   SDFFRQX2M \Rptr_reg[1]  (.SI(Rptr[0]), 
	.SE(FE_OFN24_SE), 
	.RN(R_RST), 
	.Q(Rptr[1]), 
	.D(n29), 
	.CK(R_CLK));
   SDFFRQX2M \Rptr_reg[2]  (.SI(Rptr[1]), 
	.SE(FE_OFN24_SE), 
	.RN(R_RST), 
	.Q(Rptr[2]), 
	.D(n27), 
	.CK(R_CLK));
   SDFFRQX2M \Rptr_reg[4]  (.SI(N115), 
	.SE(FE_OFN24_SE), 
	.RN(R_RST), 
	.Q(Rptr[4]), 
	.D(n31), 
	.CK(R_CLK));
   CLKINVX2M U5 (.Y(n6), 
	.A(R_RST));
   OAI2BB2X1M U6 (.Y(n25), 
	.B1(n38), 
	.B0(n7), 
	.A1N(n7), 
	.A0N(N43));
   OAI2BB2X1M U7 (.Y(n27), 
	.B1(n37), 
	.B0(n7), 
	.A1N(n7), 
	.A0N(N42));
   OAI2BB2X1M U8 (.Y(n29), 
	.B1(n36), 
	.B0(n7), 
	.A1N(n7), 
	.A0N(N41));
   NOR2BX2M U9 (.Y(\eq_41/A[1] ), 
	.B(gray_Wptr[4]), 
	.AN(n13));
   NOR2X4M U10 (.Y(Raddr[3]), 
	.B(n6), 
	.A(n38));
   NOR2X4M U11 (.Y(Raddr[0]), 
	.B(n6), 
	.A(n35));
   NOR2X4M U12 (.Y(Raddr[1]), 
	.B(n6), 
	.A(n36));
   NOR2X2M U13 (.Y(Raddr[2]), 
	.B(n6), 
	.A(n37));
   NOR2BX2M U14 (.Y(n7), 
	.B(REMPTY), 
	.AN(R_INC));
   OAI32X1M U15 (.Y(Wptr[0]), 
	.B1(n34), 
	.B0(gray_Wptr[0]), 
	.A2(n13), 
	.A1(gray_Wptr[4]), 
	.A0(n15));
   INVX2M U16 (.Y(n15), 
	.A(gray_Wptr[0]));
   INVX2M U17 (.Y(n34), 
	.A(\eq_41/A[1] ));
   XOR3XLM U18 (.Y(n13), 
	.C(gray_Wptr[2]), 
	.B(gray_Wptr[1]), 
	.A(gray_Wptr[3]));
   OAI2B2X1M U19 (.Y(n33), 
	.B1(n35), 
	.B0(n7), 
	.A1N(n7), 
	.A0(Rptr[0]));
   AO2B2X2M U20 (.Y(n31), 
	.B1(n7), 
	.B0(N44), 
	.A1N(n7), 
	.A0(Rptr[4]));
   NOR2BX2M U21 (.Y(Wptr[3]), 
	.B(gray_Wptr[4]), 
	.AN(gray_Wptr[3]));
   NOR2X2M U22 (.Y(Wptr[2]), 
	.B(n11), 
	.A(gray_Wptr[4]));
   XNOR2X2M U23 (.Y(n11), 
	.B(gray_Wptr[3]), 
	.A(gray_Wptr[2]));
   INVX2M U24 (.Y(n38), 
	.A(N115));
   INVX2M U25 (.Y(n36), 
	.A(Rptr[1]));
   INVX2M U26 (.Y(n35), 
	.A(Rptr[0]));
   OAI2BB2X1M U27 (.Y(n23), 
	.B1(n38), 
	.B0(Rptr[4]), 
	.A1N(Rptr[4]), 
	.A0N(gray_Rptr[3]));
   OAI2BB2X1M U28 (.Y(n17), 
	.B1(n3), 
	.B0(Rptr[4]), 
	.A1N(Rptr[4]), 
	.A0N(gray_Rptr[0]));
   XNOR2X2M U29 (.Y(n3), 
	.B(Rptr[1]), 
	.A(Rptr[0]));
   OAI2BB2X1M U30 (.Y(n19), 
	.B1(n4), 
	.B0(Rptr[4]), 
	.A1N(Rptr[4]), 
	.A0N(gray_Rptr[1]));
   XNOR2X2M U31 (.Y(n4), 
	.B(Rptr[2]), 
	.A(Rptr[1]));
   OAI2BB2X1M U32 (.Y(n21), 
	.B1(n5), 
	.B0(Rptr[4]), 
	.A1N(Rptr[4]), 
	.A0N(gray_Rptr[2]));
   XNOR2X2M U33 (.Y(n5), 
	.B(Rptr[2]), 
	.A(N115));
   INVX2M U44 (.Y(n37), 
	.A(Rptr[2]));
   ADDHX1M U45 (.S(N42), 
	.CO(\add_65/carry[3] ), 
	.B(\add_65/carry[2] ), 
	.A(Rptr[2]));
   ADDHX1M U46 (.S(N41), 
	.CO(\add_65/carry[2] ), 
	.B(Rptr[0]), 
	.A(Rptr[1]));
   ADDHX1M U47 (.S(N43), 
	.CO(\add_65/carry[4] ), 
	.B(\add_65/carry[3] ), 
	.A(N115));
   CLKXOR2X2M U48 (.Y(N44), 
	.B(Rptr[4]), 
	.A(\add_65/carry[4] ));
   XNOR2X1M U49 (.Y(n9), 
	.B(Wptr[2]), 
	.A(Rptr[2]));
   XNOR2X1M U50 (.Y(n8), 
	.B(Wptr[3]), 
	.A(N115));
   CLKNAND2X2M U51 (.Y(n14), 
	.B(n8), 
	.A(n9));
   CLKXOR2X2M U52 (.Y(n12), 
	.B(\eq_41/A[1] ), 
	.A(Rptr[1]));
   CLKXOR2X2M U53 (.Y(n10), 
	.B(Wptr[0]), 
	.A(Rptr[0]));
   NOR4X1M U54 (.Y(REMPTY), 
	.D(n10), 
	.C(Rptr[4]), 
	.B(n12), 
	.A(n14));
   INVX2M U3 (.Y(gray_Rptr[4]), 
	.A(HTIE_LTIEHI_NET));
endmodule

module FIFO_MEMORY_00000008_00000010_test_1 (
	WCLK, 
	WRST, 
	R_CLK, 
	R_RST, 
	wdata, 
	wclk_en, 
	rclk_en, 
	waddr, 
	raddr, 
	rdata, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN11_RST_D1_M, 
	FE_OFN12_RST_D1_M, 
	FE_OFN17_SE, 
	FE_OFN21_SE, 
	FE_OFN24_SE, 
	REF_CLK_M__L5_N2, 
	REF_CLK_M__L5_N3, 
	REF_CLK_M__L5_N4, 
	REF_CLK_M__L5_N7);
   input WCLK;
   input WRST;
   input R_CLK;
   input R_RST;
   input [7:0] wdata;
   input wclk_en;
   input rclk_en;
   input [3:0] waddr;
   input [3:0] raddr;
   output [7:0] rdata;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN11_RST_D1_M;
   input FE_OFN12_RST_D1_M;
   input FE_OFN17_SE;
   input FE_OFN21_SE;
   input FE_OFN24_SE;
   input REF_CLK_M__L5_N2;
   input REF_CLK_M__L5_N3;
   input REF_CLK_M__L5_N4;
   input REF_CLK_M__L5_N7;

   // Internal wires
   wire FE_OFN23_SE;
   wire FE_OFN13_RST_D1_M;
   wire FE_OFN9_RST_D1_M;
   wire FE_OFN7_n27;
   wire FE_OFN6_n26;
   wire FE_OFN5_n25;
   wire FE_OFN4_n24;
   wire FE_OFN3_n23;
   wire FE_OFN2_n22;
   wire FE_OFN1_n21;
   wire FE_OFN0_n3;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire \FIFO_MEM[15][7] ;
   wire \FIFO_MEM[15][6] ;
   wire \FIFO_MEM[15][5] ;
   wire \FIFO_MEM[15][4] ;
   wire \FIFO_MEM[15][3] ;
   wire \FIFO_MEM[15][2] ;
   wire \FIFO_MEM[15][1] ;
   wire \FIFO_MEM[15][0] ;
   wire \FIFO_MEM[14][7] ;
   wire \FIFO_MEM[14][6] ;
   wire \FIFO_MEM[14][5] ;
   wire \FIFO_MEM[14][4] ;
   wire \FIFO_MEM[14][3] ;
   wire \FIFO_MEM[14][2] ;
   wire \FIFO_MEM[14][1] ;
   wire \FIFO_MEM[14][0] ;
   wire \FIFO_MEM[13][7] ;
   wire \FIFO_MEM[13][6] ;
   wire \FIFO_MEM[13][5] ;
   wire \FIFO_MEM[13][4] ;
   wire \FIFO_MEM[13][3] ;
   wire \FIFO_MEM[13][2] ;
   wire \FIFO_MEM[13][1] ;
   wire \FIFO_MEM[13][0] ;
   wire \FIFO_MEM[12][7] ;
   wire \FIFO_MEM[12][6] ;
   wire \FIFO_MEM[12][5] ;
   wire \FIFO_MEM[12][4] ;
   wire \FIFO_MEM[12][3] ;
   wire \FIFO_MEM[12][2] ;
   wire \FIFO_MEM[12][1] ;
   wire \FIFO_MEM[12][0] ;
   wire \FIFO_MEM[11][7] ;
   wire \FIFO_MEM[11][6] ;
   wire \FIFO_MEM[11][5] ;
   wire \FIFO_MEM[11][4] ;
   wire \FIFO_MEM[11][3] ;
   wire \FIFO_MEM[11][2] ;
   wire \FIFO_MEM[11][1] ;
   wire \FIFO_MEM[11][0] ;
   wire \FIFO_MEM[10][7] ;
   wire \FIFO_MEM[10][6] ;
   wire \FIFO_MEM[10][5] ;
   wire \FIFO_MEM[10][4] ;
   wire \FIFO_MEM[10][3] ;
   wire \FIFO_MEM[10][2] ;
   wire \FIFO_MEM[10][1] ;
   wire \FIFO_MEM[10][0] ;
   wire \FIFO_MEM[9][7] ;
   wire \FIFO_MEM[9][6] ;
   wire \FIFO_MEM[9][5] ;
   wire \FIFO_MEM[9][4] ;
   wire \FIFO_MEM[9][3] ;
   wire \FIFO_MEM[9][2] ;
   wire \FIFO_MEM[9][1] ;
   wire \FIFO_MEM[9][0] ;
   wire \FIFO_MEM[8][7] ;
   wire \FIFO_MEM[8][6] ;
   wire \FIFO_MEM[8][5] ;
   wire \FIFO_MEM[8][4] ;
   wire \FIFO_MEM[8][3] ;
   wire \FIFO_MEM[8][2] ;
   wire \FIFO_MEM[8][1] ;
   wire \FIFO_MEM[8][0] ;
   wire \FIFO_MEM[7][7] ;
   wire \FIFO_MEM[7][6] ;
   wire \FIFO_MEM[7][5] ;
   wire \FIFO_MEM[7][4] ;
   wire \FIFO_MEM[7][3] ;
   wire \FIFO_MEM[7][2] ;
   wire \FIFO_MEM[7][1] ;
   wire \FIFO_MEM[7][0] ;
   wire \FIFO_MEM[6][7] ;
   wire \FIFO_MEM[6][6] ;
   wire \FIFO_MEM[6][5] ;
   wire \FIFO_MEM[6][4] ;
   wire \FIFO_MEM[6][3] ;
   wire \FIFO_MEM[6][2] ;
   wire \FIFO_MEM[6][1] ;
   wire \FIFO_MEM[6][0] ;
   wire \FIFO_MEM[5][7] ;
   wire \FIFO_MEM[5][6] ;
   wire \FIFO_MEM[5][5] ;
   wire \FIFO_MEM[5][4] ;
   wire \FIFO_MEM[5][3] ;
   wire \FIFO_MEM[5][2] ;
   wire \FIFO_MEM[5][1] ;
   wire \FIFO_MEM[5][0] ;
   wire \FIFO_MEM[4][7] ;
   wire \FIFO_MEM[4][6] ;
   wire \FIFO_MEM[4][5] ;
   wire \FIFO_MEM[4][4] ;
   wire \FIFO_MEM[4][3] ;
   wire \FIFO_MEM[4][2] ;
   wire \FIFO_MEM[4][1] ;
   wire \FIFO_MEM[4][0] ;
   wire \FIFO_MEM[3][7] ;
   wire \FIFO_MEM[3][6] ;
   wire \FIFO_MEM[3][5] ;
   wire \FIFO_MEM[3][4] ;
   wire \FIFO_MEM[3][3] ;
   wire \FIFO_MEM[3][2] ;
   wire \FIFO_MEM[3][1] ;
   wire \FIFO_MEM[3][0] ;
   wire \FIFO_MEM[2][7] ;
   wire \FIFO_MEM[2][6] ;
   wire \FIFO_MEM[2][5] ;
   wire \FIFO_MEM[2][4] ;
   wire \FIFO_MEM[2][3] ;
   wire \FIFO_MEM[2][2] ;
   wire \FIFO_MEM[2][1] ;
   wire \FIFO_MEM[2][0] ;
   wire \FIFO_MEM[1][7] ;
   wire \FIFO_MEM[1][6] ;
   wire \FIFO_MEM[1][5] ;
   wire \FIFO_MEM[1][4] ;
   wire \FIFO_MEM[1][3] ;
   wire \FIFO_MEM[1][2] ;
   wire \FIFO_MEM[1][1] ;
   wire \FIFO_MEM[1][0] ;
   wire \FIFO_MEM[0][7] ;
   wire \FIFO_MEM[0][6] ;
   wire \FIFO_MEM[0][5] ;
   wire \FIFO_MEM[0][4] ;
   wire \FIFO_MEM[0][3] ;
   wire \FIFO_MEM[0][2] ;
   wire \FIFO_MEM[0][1] ;
   wire \FIFO_MEM[0][0] ;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N57;
   wire N58;
   wire N59;
   wire N60;
   wire N61;
   wire N62;
   wire N63;
   wire N64;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n35;
   wire n36;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n47;
   wire n49;
   wire n51;
   wire n53;
   wire n55;
   wire n57;
   wire n59;
   wire n61;
   wire n63;
   wire n65;
   wire n67;
   wire n69;
   wire n71;
   wire n73;
   wire n75;
   wire n77;
   wire n80;
   wire n82;
   wire n84;
   wire n86;
   wire n88;
   wire n90;
   wire n92;
   wire n94;
   wire n96;
   wire n98;
   wire n100;
   wire n102;
   wire n104;
   wire n106;
   wire n108;
   wire n110;
   wire n113;
   wire n115;
   wire n117;
   wire n119;
   wire n121;
   wire n123;
   wire n125;
   wire n127;
   wire n129;
   wire n131;
   wire n133;
   wire n135;
   wire n137;
   wire n139;
   wire n141;
   wire n143;
   wire n146;
   wire n148;
   wire n150;
   wire n152;
   wire n154;
   wire n156;
   wire n158;
   wire n160;
   wire n162;
   wire n164;
   wire n166;
   wire n168;
   wire n170;
   wire n172;
   wire n174;
   wire n176;
   wire n179;
   wire n181;
   wire n183;
   wire n185;
   wire n187;
   wire n189;
   wire n191;
   wire n193;
   wire n195;
   wire n197;
   wire n199;
   wire n201;
   wire n203;
   wire n205;
   wire n207;
   wire n209;
   wire n212;
   wire n214;
   wire n216;
   wire n218;
   wire n220;
   wire n222;
   wire n224;
   wire n226;
   wire n228;
   wire n230;
   wire n232;
   wire n234;
   wire n236;
   wire n238;
   wire n240;
   wire n242;
   wire n245;
   wire n247;
   wire n249;
   wire n251;
   wire n253;
   wire n255;
   wire n257;
   wire n259;
   wire n261;
   wire n263;
   wire n265;
   wire n267;
   wire n269;
   wire n271;
   wire n273;
   wire n275;
   wire n278;
   wire n280;
   wire n282;
   wire n284;
   wire n286;
   wire n288;
   wire n290;
   wire n292;
   wire n294;
   wire n296;
   wire n298;
   wire n300;
   wire n302;
   wire n304;
   wire n306;
   wire n308;
   wire n34;
   wire n37;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n350;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n387;
   wire n388;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n419;
   wire n420;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire [7:0] out_next;

   assign N11 = raddr[0] ;
   assign N12 = raddr[1] ;
   assign N13 = raddr[2] ;
   assign N14 = raddr[3] ;
   assign N15 = waddr[0] ;
   assign N16 = waddr[1] ;
   assign N17 = waddr[2] ;
   assign N18 = waddr[3] ;
   assign test_so1 = \FIFO_MEM[9][6]  ;

   CLKBUFX6M FE_OFC23_SE (.Y(FE_OFN23_SE), 
	.A(FE_OFN17_SE));
   BUFX6M FE_OFC13_RST_D1_M (.Y(FE_OFN13_RST_D1_M), 
	.A(FE_OFN9_RST_D1_M));
   BUFX5M FE_OFC9_RST_D1_M (.Y(FE_OFN9_RST_D1_M), 
	.A(WRST));
   BUFX2M FE_OFC7_n27 (.Y(FE_OFN7_n27), 
	.A(n27));
   BUFX2M FE_OFC6_n26 (.Y(FE_OFN6_n26), 
	.A(n26));
   BUFX2M FE_OFC5_n25 (.Y(FE_OFN5_n25), 
	.A(n25));
   BUFX2M FE_OFC4_n24 (.Y(FE_OFN4_n24), 
	.A(n24));
   BUFX2M FE_OFC3_n23 (.Y(FE_OFN3_n23), 
	.A(n23));
   BUFX2M FE_OFC2_n22 (.Y(FE_OFN2_n22), 
	.A(n22));
   BUFX2M FE_OFC1_n21 (.Y(FE_OFN1_n21), 
	.A(n21));
   BUFX2M FE_OFC0_n3 (.Y(FE_OFN0_n3), 
	.A(n3));
   SDFFRQX2M \out_next_reg[7]  (.SI(out_next[6]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(out_next[7]), 
	.D(N57), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \out_next_reg[6]  (.SI(out_next[5]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(out_next[6]), 
	.D(N58), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \out_next_reg[5]  (.SI(out_next[4]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(out_next[5]), 
	.D(N59), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \out_next_reg[4]  (.SI(out_next[3]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(out_next[4]), 
	.D(N60), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \out_next_reg[3]  (.SI(out_next[2]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(out_next[3]), 
	.D(N61), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \out_next_reg[2]  (.SI(out_next[1]), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(out_next[2]), 
	.D(N62), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \out_next_reg[1]  (.SI(out_next[0]), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(out_next[1]), 
	.D(N63), 
	.CK(WCLK));
   SDFFRQX2M \out_next_reg[0]  (.SI(\FIFO_MEM[15][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(out_next[0]), 
	.D(N64), 
	.CK(REF_CLK_M__L5_N4));
   SEDFFX2M \read_next_reg[7]  (.SI(n422), 
	.SE(FE_OFN24_SE), 
	.QN(n45), 
	.Q(test_so2), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[7]), 
	.CK(REF_CLK_M__L5_N4));
   SEDFFX2M \read_next_reg[6]  (.SI(n423), 
	.SE(FE_OFN24_SE), 
	.QN(n44), 
	.Q(n422), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[6]), 
	.CK(REF_CLK_M__L5_N4));
   SEDFFX2M \read_next_reg[4]  (.SI(n425), 
	.SE(FE_OFN24_SE), 
	.QN(n42), 
	.Q(n424), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[4]), 
	.CK(REF_CLK_M__L5_N4));
   SEDFFX2M \read_next_reg[3]  (.SI(n426), 
	.SE(FE_OFN24_SE), 
	.QN(n41), 
	.Q(n425), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[3]), 
	.CK(REF_CLK_M__L5_N4));
   SEDFFX2M \read_next_reg[2]  (.SI(n427), 
	.SE(FE_OFN24_SE), 
	.QN(n40), 
	.Q(n426), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[2]), 
	.CK(REF_CLK_M__L5_N4));
   SEDFFX2M \read_next_reg[1]  (.SI(n428), 
	.SE(FE_OFN24_SE), 
	.QN(n39), 
	.Q(n427), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[1]), 
	.CK(REF_CLK_M__L5_N4));
   SEDFFX2M \read_next_reg[0]  (.SI(out_next[7]), 
	.SE(FE_OFN24_SE), 
	.QN(n38), 
	.Q(n428), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[0]), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[13][7]  (.SI(\FIFO_MEM[13][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][7] ), 
	.D(n304), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][7]  (.SI(test_si2), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[9][7] ), 
	.D(n296), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[5][7]  (.SI(\FIFO_MEM[5][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][7] ), 
	.D(n288), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[1][7]  (.SI(\FIFO_MEM[1][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[1][7] ), 
	.D(n280), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[13][6]  (.SI(\FIFO_MEM[13][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][6] ), 
	.D(n271), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][6]  (.SI(\FIFO_MEM[9][5] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[9][6] ), 
	.D(n263), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[5][6]  (.SI(\FIFO_MEM[5][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][6] ), 
	.D(n255), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[1][6]  (.SI(\FIFO_MEM[1][5] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[1][6] ), 
	.D(n247), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[13][5]  (.SI(\FIFO_MEM[13][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][5] ), 
	.D(n238), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][5]  (.SI(\FIFO_MEM[9][4] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[9][5] ), 
	.D(n230), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[5][5]  (.SI(\FIFO_MEM[5][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][5] ), 
	.D(n222), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[1][5]  (.SI(\FIFO_MEM[1][4] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[1][5] ), 
	.D(n214), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[13][4]  (.SI(\FIFO_MEM[13][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][4] ), 
	.D(n205), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][4]  (.SI(\FIFO_MEM[9][3] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[9][4] ), 
	.D(n197), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[5][4]  (.SI(\FIFO_MEM[5][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][4] ), 
	.D(n189), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[1][4]  (.SI(\FIFO_MEM[1][3] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[1][4] ), 
	.D(n181), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[13][3]  (.SI(\FIFO_MEM[13][2] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][3] ), 
	.D(n172), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][3]  (.SI(\FIFO_MEM[9][2] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[9][3] ), 
	.D(n164), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[5][3]  (.SI(\FIFO_MEM[5][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][3] ), 
	.D(n156), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[1][3]  (.SI(\FIFO_MEM[1][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[1][3] ), 
	.D(n148), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[13][2]  (.SI(\FIFO_MEM[13][1] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][2] ), 
	.D(n139), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][2]  (.SI(\FIFO_MEM[9][1] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[9][2] ), 
	.D(n131), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[5][2]  (.SI(\FIFO_MEM[5][1] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][2] ), 
	.D(n123), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[1][2]  (.SI(\FIFO_MEM[1][1] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[1][2] ), 
	.D(n115), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[13][1]  (.SI(\FIFO_MEM[13][0] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][1] ), 
	.D(n106), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][1]  (.SI(\FIFO_MEM[9][0] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[9][1] ), 
	.D(n98), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[5][1]  (.SI(\FIFO_MEM[5][0] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][1] ), 
	.D(n90), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[1][1]  (.SI(\FIFO_MEM[1][0] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[1][1] ), 
	.D(n82), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[13][0]  (.SI(\FIFO_MEM[12][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[13][0] ), 
	.D(n73), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[9][0]  (.SI(\FIFO_MEM[8][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[9][0] ), 
	.D(n65), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[5][0]  (.SI(\FIFO_MEM[4][7] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[5][0] ), 
	.D(n57), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[1][0]  (.SI(\FIFO_MEM[0][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[1][0] ), 
	.D(n49), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[15][7]  (.SI(\FIFO_MEM[15][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][7] ), 
	.D(n308), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][7]  (.SI(\FIFO_MEM[11][6] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[11][7] ), 
	.D(n300), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[7][7]  (.SI(\FIFO_MEM[7][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[7][7] ), 
	.D(n292), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[3][7]  (.SI(\FIFO_MEM[3][6] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[3][7] ), 
	.D(n284), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[15][6]  (.SI(\FIFO_MEM[15][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][6] ), 
	.D(n275), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][6]  (.SI(\FIFO_MEM[11][5] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[11][6] ), 
	.D(n267), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[7][6]  (.SI(\FIFO_MEM[7][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[7][6] ), 
	.D(n259), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[3][6]  (.SI(\FIFO_MEM[3][5] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[3][6] ), 
	.D(n251), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[15][5]  (.SI(\FIFO_MEM[15][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][5] ), 
	.D(n242), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][5]  (.SI(\FIFO_MEM[11][4] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[11][5] ), 
	.D(n234), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[7][5]  (.SI(\FIFO_MEM[7][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[7][5] ), 
	.D(n226), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[3][5]  (.SI(\FIFO_MEM[3][4] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[3][5] ), 
	.D(n218), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[15][4]  (.SI(\FIFO_MEM[15][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][4] ), 
	.D(n209), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][4]  (.SI(\FIFO_MEM[11][3] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[11][4] ), 
	.D(n201), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[7][4]  (.SI(\FIFO_MEM[7][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[7][4] ), 
	.D(n193), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[3][4]  (.SI(\FIFO_MEM[3][3] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\FIFO_MEM[3][4] ), 
	.D(n185), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[15][3]  (.SI(\FIFO_MEM[15][2] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][3] ), 
	.D(n176), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][3]  (.SI(\FIFO_MEM[11][2] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[11][3] ), 
	.D(n168), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[7][3]  (.SI(\FIFO_MEM[7][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[7][3] ), 
	.D(n160), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[3][3]  (.SI(\FIFO_MEM[3][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[3][3] ), 
	.D(n152), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[15][2]  (.SI(\FIFO_MEM[15][1] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][2] ), 
	.D(n143), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][2]  (.SI(\FIFO_MEM[11][1] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[11][2] ), 
	.D(n135), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[7][2]  (.SI(\FIFO_MEM[7][1] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[7][2] ), 
	.D(n127), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[3][2]  (.SI(\FIFO_MEM[3][1] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[3][2] ), 
	.D(n119), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[15][1]  (.SI(\FIFO_MEM[15][0] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][1] ), 
	.D(n110), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][1]  (.SI(\FIFO_MEM[11][0] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[11][1] ), 
	.D(n102), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[7][1]  (.SI(\FIFO_MEM[7][0] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[7][1] ), 
	.D(n94), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[3][1]  (.SI(\FIFO_MEM[3][0] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[3][1] ), 
	.D(n86), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[15][0]  (.SI(\FIFO_MEM[14][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[15][0] ), 
	.D(n77), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[11][0]  (.SI(\FIFO_MEM[10][7] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[11][0] ), 
	.D(n69), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[7][0]  (.SI(\FIFO_MEM[6][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[7][0] ), 
	.D(n61), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[3][0]  (.SI(\FIFO_MEM[2][7] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[3][0] ), 
	.D(n53), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[14][7]  (.SI(\FIFO_MEM[14][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][7] ), 
	.D(n306), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][7]  (.SI(\FIFO_MEM[10][6] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[10][7] ), 
	.D(n298), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][7]  (.SI(\FIFO_MEM[6][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][7] ), 
	.D(n290), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][7]  (.SI(\FIFO_MEM[2][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[2][7] ), 
	.D(n282), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[14][6]  (.SI(\FIFO_MEM[14][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][6] ), 
	.D(n273), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][6]  (.SI(\FIFO_MEM[10][5] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[10][6] ), 
	.D(n265), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][6]  (.SI(\FIFO_MEM[6][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][6] ), 
	.D(n257), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][6]  (.SI(\FIFO_MEM[2][5] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[2][6] ), 
	.D(n249), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[14][5]  (.SI(\FIFO_MEM[14][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][5] ), 
	.D(n240), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][5]  (.SI(\FIFO_MEM[10][4] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[10][5] ), 
	.D(n232), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][5]  (.SI(\FIFO_MEM[6][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][5] ), 
	.D(n224), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][5]  (.SI(\FIFO_MEM[2][4] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[2][5] ), 
	.D(n216), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[14][4]  (.SI(\FIFO_MEM[14][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][4] ), 
	.D(n207), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][4]  (.SI(\FIFO_MEM[10][3] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[10][4] ), 
	.D(n199), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][4]  (.SI(\FIFO_MEM[6][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][4] ), 
	.D(n191), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][4]  (.SI(\FIFO_MEM[2][3] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[2][4] ), 
	.D(n183), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[14][3]  (.SI(\FIFO_MEM[14][2] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][3] ), 
	.D(n174), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][3]  (.SI(\FIFO_MEM[10][2] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[10][3] ), 
	.D(n166), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][3]  (.SI(\FIFO_MEM[6][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][3] ), 
	.D(n158), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][3]  (.SI(\FIFO_MEM[2][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[2][3] ), 
	.D(n150), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[14][2]  (.SI(\FIFO_MEM[14][1] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][2] ), 
	.D(n141), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][2]  (.SI(\FIFO_MEM[10][1] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[10][2] ), 
	.D(n133), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][2]  (.SI(\FIFO_MEM[6][1] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][2] ), 
	.D(n125), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][2]  (.SI(\FIFO_MEM[2][1] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[2][2] ), 
	.D(n117), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[14][1]  (.SI(\FIFO_MEM[14][0] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][1] ), 
	.D(n108), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][1]  (.SI(\FIFO_MEM[10][0] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[10][1] ), 
	.D(n100), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][1]  (.SI(\FIFO_MEM[6][0] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][1] ), 
	.D(n92), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][1]  (.SI(\FIFO_MEM[2][0] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[2][1] ), 
	.D(n84), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[14][0]  (.SI(\FIFO_MEM[13][7] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[14][0] ), 
	.D(n75), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[10][0]  (.SI(\FIFO_MEM[9][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[10][0] ), 
	.D(n67), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[6][0]  (.SI(\FIFO_MEM[5][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[6][0] ), 
	.D(n59), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[2][0]  (.SI(\FIFO_MEM[1][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[2][0] ), 
	.D(n51), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[12][7]  (.SI(\FIFO_MEM[12][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][7] ), 
	.D(n302), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][7]  (.SI(\FIFO_MEM[8][6] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[8][7] ), 
	.D(n294), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[4][7]  (.SI(\FIFO_MEM[4][6] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[4][7] ), 
	.D(n286), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][7]  (.SI(\FIFO_MEM[0][6] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[0][7] ), 
	.D(n278), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[12][6]  (.SI(\FIFO_MEM[12][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][6] ), 
	.D(n269), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][6]  (.SI(\FIFO_MEM[8][5] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[8][6] ), 
	.D(n261), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[4][6]  (.SI(\FIFO_MEM[4][5] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[4][6] ), 
	.D(n253), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][6]  (.SI(\FIFO_MEM[0][5] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[0][6] ), 
	.D(n245), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[12][5]  (.SI(\FIFO_MEM[12][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][5] ), 
	.D(n236), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][5]  (.SI(\FIFO_MEM[8][4] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[8][5] ), 
	.D(n228), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[4][5]  (.SI(\FIFO_MEM[4][4] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[4][5] ), 
	.D(n220), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][5]  (.SI(\FIFO_MEM[0][4] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[0][5] ), 
	.D(n212), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[12][4]  (.SI(\FIFO_MEM[12][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][4] ), 
	.D(n203), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][4]  (.SI(\FIFO_MEM[8][3] ), 
	.SE(FE_OFN17_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[8][4] ), 
	.D(n195), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[4][4]  (.SI(\FIFO_MEM[4][3] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[4][4] ), 
	.D(n187), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][4]  (.SI(\FIFO_MEM[0][3] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\FIFO_MEM[0][4] ), 
	.D(n179), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[12][3]  (.SI(\FIFO_MEM[12][2] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][3] ), 
	.D(n170), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][3]  (.SI(\FIFO_MEM[8][2] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[8][3] ), 
	.D(n162), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[4][3]  (.SI(\FIFO_MEM[4][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[4][3] ), 
	.D(n154), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][3]  (.SI(\FIFO_MEM[0][2] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\FIFO_MEM[0][3] ), 
	.D(n146), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[12][2]  (.SI(\FIFO_MEM[12][1] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][2] ), 
	.D(n137), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][2]  (.SI(\FIFO_MEM[8][1] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[8][2] ), 
	.D(n129), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[4][2]  (.SI(\FIFO_MEM[4][1] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[4][2] ), 
	.D(n121), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][2]  (.SI(\FIFO_MEM[0][1] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[0][2] ), 
	.D(n113), 
	.CK(WCLK));
   SDFFRQX2M \FIFO_MEM_reg[12][1]  (.SI(\FIFO_MEM[12][0] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][1] ), 
	.D(n104), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][1]  (.SI(\FIFO_MEM[8][0] ), 
	.SE(FE_OFN24_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[8][1] ), 
	.D(n96), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[4][1]  (.SI(\FIFO_MEM[4][0] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[4][1] ), 
	.D(n88), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][1]  (.SI(\FIFO_MEM[0][0] ), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\FIFO_MEM[0][1] ), 
	.D(n80), 
	.CK(REF_CLK_M__L5_N2));
   SDFFRQX2M \FIFO_MEM_reg[12][0]  (.SI(\FIFO_MEM[11][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN13_RST_D1_M), 
	.Q(\FIFO_MEM[12][0] ), 
	.D(n71), 
	.CK(REF_CLK_M__L5_N7));
   SDFFRQX2M \FIFO_MEM_reg[8][0]  (.SI(\FIFO_MEM[7][7] ), 
	.SE(FE_OFN23_SE), 
	.RN(FE_OFN9_RST_D1_M), 
	.Q(\FIFO_MEM[8][0] ), 
	.D(n63), 
	.CK(REF_CLK_M__L5_N4));
   SDFFRQX2M \FIFO_MEM_reg[4][0]  (.SI(\FIFO_MEM[3][7] ), 
	.SE(FE_OFN21_SE), 
	.RN(FE_OFN12_RST_D1_M), 
	.Q(\FIFO_MEM[4][0] ), 
	.D(n55), 
	.CK(REF_CLK_M__L5_N3));
   SDFFRQX2M \FIFO_MEM_reg[0][0]  (.SI(test_si1), 
	.SE(test_se), 
	.RN(FE_OFN11_RST_D1_M), 
	.Q(\FIFO_MEM[0][0] ), 
	.D(n47), 
	.CK(REF_CLK_M__L5_N2));
   SEDFFX1M \read_next_reg[5]  (.SI(n424), 
	.SE(FE_OFN24_SE), 
	.QN(n43), 
	.Q(n423), 
	.E(FE_OFN12_RST_D1_M), 
	.D(rdata[5]), 
	.CK(REF_CLK_M__L5_N4));
   NOR2X2M U4 (.Y(n30), 
	.B(n399), 
	.A(n398));
   NOR2X2M U5 (.Y(n29), 
	.B(n399), 
	.A(N15));
   INVX4M U6 (.Y(n387), 
	.A(n398));
   INVX4M U7 (.Y(n388), 
	.A(n398));
   INVX3M U22 (.Y(n350), 
	.A(n348));
   INVX2M U27 (.Y(n419), 
	.A(wclk_en));
   NOR2X2M U28 (.Y(n33), 
	.B(N18), 
	.A(n420));
   NAND2X2M U29 (.Y(n10), 
	.B(n31), 
	.A(n33));
   NAND2X2M U30 (.Y(n11), 
	.B(n32), 
	.A(n33));
   NAND2X2M U31 (.Y(n14), 
	.B(n31), 
	.A(n35));
   NAND2X2M U32 (.Y(n15), 
	.B(n32), 
	.A(n35));
   NAND2X2M U33 (.Y(n18), 
	.B(n31), 
	.A(n36));
   NAND2X2M U34 (.Y(n19), 
	.B(n32), 
	.A(n36));
   NAND2X2M U35 (.Y(n8), 
	.B(n29), 
	.A(n33));
   NAND2X2M U36 (.Y(n9), 
	.B(n30), 
	.A(n33));
   NAND2X2M U37 (.Y(n12), 
	.B(n29), 
	.A(n35));
   NAND2X2M U38 (.Y(n13), 
	.B(n30), 
	.A(n35));
   NAND2X2M U39 (.Y(n16), 
	.B(n29), 
	.A(n36));
   NAND2X2M U40 (.Y(n17), 
	.B(n30), 
	.A(n36));
   AND2X2M U41 (.Y(n35), 
	.B(n420), 
	.A(N18));
   AND2X2M U42 (.Y(n36), 
	.B(N17), 
	.A(N18));
   INVX2M U43 (.Y(n420), 
	.A(N17));
   NOR2X2M U46 (.Y(n28), 
	.B(N18), 
	.A(N17));
   NAND2X2M U47 (.Y(n5), 
	.B(n28), 
	.A(n30));
   NAND2X2M U48 (.Y(n6), 
	.B(n28), 
	.A(n31));
   NAND2X2M U49 (.Y(n7), 
	.B(n28), 
	.A(n32));
   NAND2X2M U50 (.Y(n4), 
	.B(n29), 
	.A(n28));
   NAND2BX2M U53 (.Y(n1), 
	.B(R_RST), 
	.AN(rclk_en));
   AND2X2M U54 (.Y(n2), 
	.B(R_RST), 
	.A(rclk_en));
   INVX2M U55 (.Y(n398), 
	.A(N15));
   BUFX6M U57 (.Y(n397), 
	.A(N11));
   INVX2M U58 (.Y(n348), 
	.A(N12));
   AND2X2M U59 (.Y(n31), 
	.B(n398), 
	.A(n399));
   AND2X2M U60 (.Y(n32), 
	.B(N15), 
	.A(n399));
   OAI2BB2X1M U61 (.Y(rdata[2]), 
	.B1(n40), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N53));
   MX4X1M U62 (.Y(N53), 
	.S1(N13), 
	.S0(N14), 
	.D(n324), 
	.C(n326), 
	.B(n325), 
	.A(n327));
   MX4X1M U63 (.Y(n327), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[3][2] ), 
	.C(\FIFO_MEM[2][2] ), 
	.B(\FIFO_MEM[1][2] ), 
	.A(\FIFO_MEM[0][2] ));
   MX4X1M U64 (.Y(n325), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[11][2] ), 
	.C(\FIFO_MEM[10][2] ), 
	.B(\FIFO_MEM[9][2] ), 
	.A(\FIFO_MEM[8][2] ));
   OAI2BB2X1M U65 (.Y(rdata[6]), 
	.B1(n44), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N49));
   MX4X1M U66 (.Y(N49), 
	.S1(N13), 
	.S0(N14), 
	.D(n340), 
	.C(n342), 
	.B(n341), 
	.A(n343));
   MX4X1M U67 (.Y(n343), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[3][6] ), 
	.C(\FIFO_MEM[2][6] ), 
	.B(\FIFO_MEM[1][6] ), 
	.A(\FIFO_MEM[0][6] ));
   MX4X1M U68 (.Y(n341), 
	.S1(N12), 
	.S0(N11), 
	.D(\FIFO_MEM[11][6] ), 
	.C(\FIFO_MEM[10][6] ), 
	.B(\FIFO_MEM[9][6] ), 
	.A(\FIFO_MEM[8][6] ));
   OAI2BB2X1M U69 (.Y(rdata[3]), 
	.B1(n41), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N52));
   MX4X1M U70 (.Y(N52), 
	.S1(N13), 
	.S0(N14), 
	.D(n328), 
	.C(n330), 
	.B(n329), 
	.A(n331));
   MX4X1M U71 (.Y(n331), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[3][3] ), 
	.C(\FIFO_MEM[2][3] ), 
	.B(\FIFO_MEM[1][3] ), 
	.A(\FIFO_MEM[0][3] ));
   MX4X1M U72 (.Y(n329), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[11][3] ), 
	.C(\FIFO_MEM[10][3] ), 
	.B(\FIFO_MEM[9][3] ), 
	.A(\FIFO_MEM[8][3] ));
   OAI2BB2X1M U73 (.Y(rdata[7]), 
	.B1(n45), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N48));
   MX4X1M U74 (.Y(N48), 
	.S1(N13), 
	.S0(N14), 
	.D(n344), 
	.C(n346), 
	.B(n345), 
	.A(n347));
   MX4X1M U75 (.Y(n347), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[3][7] ), 
	.C(\FIFO_MEM[2][7] ), 
	.B(\FIFO_MEM[1][7] ), 
	.A(\FIFO_MEM[0][7] ));
   MX4X1M U76 (.Y(n345), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[11][7] ), 
	.C(\FIFO_MEM[10][7] ), 
	.B(\FIFO_MEM[9][7] ), 
	.A(\FIFO_MEM[8][7] ));
   OAI2BB2X1M U77 (.Y(rdata[0]), 
	.B1(n38), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N55));
   MX4X1M U78 (.Y(N55), 
	.S1(N13), 
	.S0(N14), 
	.D(n34), 
	.C(n318), 
	.B(n37), 
	.A(n319));
   MX4X1M U79 (.Y(n319), 
	.S1(N12), 
	.S0(N11), 
	.D(\FIFO_MEM[3][0] ), 
	.C(\FIFO_MEM[2][0] ), 
	.B(\FIFO_MEM[1][0] ), 
	.A(\FIFO_MEM[0][0] ));
   MX4X1M U80 (.Y(n37), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[11][0] ), 
	.C(\FIFO_MEM[10][0] ), 
	.B(\FIFO_MEM[9][0] ), 
	.A(\FIFO_MEM[8][0] ));
   OAI2BB2X1M U81 (.Y(rdata[4]), 
	.B1(n42), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N51));
   MX4X1M U82 (.Y(N51), 
	.S1(N13), 
	.S0(N14), 
	.D(n332), 
	.C(n334), 
	.B(n333), 
	.A(n335));
   MX4X1M U83 (.Y(n335), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[3][4] ), 
	.C(\FIFO_MEM[2][4] ), 
	.B(\FIFO_MEM[1][4] ), 
	.A(\FIFO_MEM[0][4] ));
   MX4X1M U84 (.Y(n333), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[11][4] ), 
	.C(\FIFO_MEM[10][4] ), 
	.B(\FIFO_MEM[9][4] ), 
	.A(\FIFO_MEM[8][4] ));
   OAI2BB2X1M U85 (.Y(rdata[1]), 
	.B1(n39), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N54));
   MX4X1M U86 (.Y(N54), 
	.S1(N13), 
	.S0(N14), 
	.D(n320), 
	.C(n322), 
	.B(n321), 
	.A(n323));
   MX4X1M U87 (.Y(n321), 
	.S1(N12), 
	.S0(N11), 
	.D(\FIFO_MEM[11][1] ), 
	.C(\FIFO_MEM[10][1] ), 
	.B(\FIFO_MEM[9][1] ), 
	.A(\FIFO_MEM[8][1] ));
   MX4X1M U88 (.Y(n320), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[15][1] ), 
	.C(\FIFO_MEM[14][1] ), 
	.B(\FIFO_MEM[13][1] ), 
	.A(\FIFO_MEM[12][1] ));
   OAI2BB2X1M U89 (.Y(rdata[5]), 
	.B1(n43), 
	.B0(n1), 
	.A1N(n2), 
	.A0N(N50));
   MX4X1M U90 (.Y(N50), 
	.S1(N13), 
	.S0(N14), 
	.D(n336), 
	.C(n338), 
	.B(n337), 
	.A(n339));
   MX4X1M U91 (.Y(n339), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[3][5] ), 
	.C(\FIFO_MEM[2][5] ), 
	.B(\FIFO_MEM[1][5] ), 
	.A(\FIFO_MEM[0][5] ));
   MX4X1M U92 (.Y(n337), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[11][5] ), 
	.C(\FIFO_MEM[10][5] ), 
	.B(\FIFO_MEM[9][5] ), 
	.A(\FIFO_MEM[8][5] ));
   AOI22X1M U94 (.Y(n3), 
	.B1(n419), 
	.B0(out_next[0]), 
	.A1(wclk_en), 
	.A0(wdata[0]));
   AOI22X1M U96 (.Y(n21), 
	.B1(n419), 
	.B0(out_next[1]), 
	.A1(wclk_en), 
	.A0(wdata[1]));
   AOI22X1M U98 (.Y(n22), 
	.B1(n419), 
	.B0(out_next[2]), 
	.A1(wclk_en), 
	.A0(wdata[2]));
   AOI22X1M U100 (.Y(n23), 
	.B1(n419), 
	.B0(out_next[3]), 
	.A1(wclk_en), 
	.A0(wdata[3]));
   AOI22X1M U102 (.Y(n24), 
	.B1(n419), 
	.B0(out_next[4]), 
	.A1(wclk_en), 
	.A0(wdata[4]));
   AOI22X1M U104 (.Y(n25), 
	.B1(n419), 
	.B0(out_next[5]), 
	.A1(wclk_en), 
	.A0(wdata[5]));
   AOI22X1M U106 (.Y(n26), 
	.B1(n419), 
	.B0(out_next[6]), 
	.A1(wclk_en), 
	.A0(wdata[6]));
   AOI22X1M U108 (.Y(n27), 
	.B1(n419), 
	.B0(out_next[7]), 
	.A1(wclk_en), 
	.A0(wdata[7]));
   OAI2BB2X1M U109 (.Y(n47), 
	.B1(n4), 
	.B0(FE_OFN0_n3), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][0] ));
   OAI2BB2X1M U110 (.Y(n49), 
	.B1(n5), 
	.B0(FE_OFN0_n3), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][0] ));
   OAI2BB2X1M U111 (.Y(n80), 
	.B1(n4), 
	.B0(FE_OFN1_n21), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][1] ));
   OAI2BB2X1M U112 (.Y(n82), 
	.B1(n5), 
	.B0(FE_OFN1_n21), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][1] ));
   OAI2BB2X1M U113 (.Y(n113), 
	.B1(n4), 
	.B0(FE_OFN2_n22), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][2] ));
   OAI2BB2X1M U114 (.Y(n115), 
	.B1(n5), 
	.B0(FE_OFN2_n22), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][2] ));
   OAI2BB2X1M U115 (.Y(n146), 
	.B1(n4), 
	.B0(FE_OFN3_n23), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][3] ));
   OAI2BB2X1M U116 (.Y(n148), 
	.B1(n5), 
	.B0(FE_OFN3_n23), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][3] ));
   OAI2BB2X1M U117 (.Y(n179), 
	.B1(n4), 
	.B0(FE_OFN4_n24), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][4] ));
   OAI2BB2X1M U118 (.Y(n181), 
	.B1(n5), 
	.B0(FE_OFN4_n24), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][4] ));
   OAI2BB2X1M U119 (.Y(n212), 
	.B1(n4), 
	.B0(FE_OFN5_n25), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][5] ));
   OAI2BB2X1M U120 (.Y(n214), 
	.B1(n5), 
	.B0(FE_OFN5_n25), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][5] ));
   OAI2BB2X1M U121 (.Y(n245), 
	.B1(n4), 
	.B0(FE_OFN6_n26), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][6] ));
   OAI2BB2X1M U122 (.Y(n247), 
	.B1(n5), 
	.B0(FE_OFN6_n26), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][6] ));
   OAI2BB2X1M U123 (.Y(n278), 
	.B1(n4), 
	.B0(FE_OFN7_n27), 
	.A1N(n4), 
	.A0N(\FIFO_MEM[0][7] ));
   OAI2BB2X1M U124 (.Y(n280), 
	.B1(n5), 
	.B0(FE_OFN7_n27), 
	.A1N(n5), 
	.A0N(\FIFO_MEM[1][7] ));
   OAI2BB2X1M U125 (.Y(n55), 
	.B1(n8), 
	.B0(FE_OFN0_n3), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][0] ));
   OAI2BB2X1M U126 (.Y(n57), 
	.B1(n9), 
	.B0(FE_OFN0_n3), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][0] ));
   OAI2BB2X1M U127 (.Y(n59), 
	.B1(n10), 
	.B0(FE_OFN0_n3), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][0] ));
   OAI2BB2X1M U128 (.Y(n61), 
	.B1(n11), 
	.B0(FE_OFN0_n3), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][0] ));
   OAI2BB2X1M U129 (.Y(n88), 
	.B1(n8), 
	.B0(FE_OFN1_n21), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][1] ));
   OAI2BB2X1M U130 (.Y(n90), 
	.B1(n9), 
	.B0(FE_OFN1_n21), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][1] ));
   OAI2BB2X1M U131 (.Y(n92), 
	.B1(n10), 
	.B0(FE_OFN1_n21), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][1] ));
   OAI2BB2X1M U132 (.Y(n94), 
	.B1(n11), 
	.B0(FE_OFN1_n21), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][1] ));
   OAI2BB2X1M U133 (.Y(n121), 
	.B1(n8), 
	.B0(FE_OFN2_n22), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][2] ));
   OAI2BB2X1M U134 (.Y(n123), 
	.B1(n9), 
	.B0(FE_OFN2_n22), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][2] ));
   OAI2BB2X1M U135 (.Y(n125), 
	.B1(n10), 
	.B0(FE_OFN2_n22), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][2] ));
   OAI2BB2X1M U136 (.Y(n127), 
	.B1(n11), 
	.B0(FE_OFN2_n22), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][2] ));
   OAI2BB2X1M U137 (.Y(n154), 
	.B1(n8), 
	.B0(FE_OFN3_n23), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][3] ));
   OAI2BB2X1M U138 (.Y(n156), 
	.B1(n9), 
	.B0(FE_OFN3_n23), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][3] ));
   OAI2BB2X1M U139 (.Y(n158), 
	.B1(n10), 
	.B0(FE_OFN3_n23), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][3] ));
   OAI2BB2X1M U140 (.Y(n160), 
	.B1(n11), 
	.B0(FE_OFN3_n23), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][3] ));
   OAI2BB2X1M U141 (.Y(n187), 
	.B1(n8), 
	.B0(FE_OFN4_n24), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][4] ));
   OAI2BB2X1M U142 (.Y(n189), 
	.B1(n9), 
	.B0(FE_OFN4_n24), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][4] ));
   OAI2BB2X1M U143 (.Y(n191), 
	.B1(n10), 
	.B0(FE_OFN4_n24), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][4] ));
   OAI2BB2X1M U144 (.Y(n193), 
	.B1(n11), 
	.B0(FE_OFN4_n24), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][4] ));
   OAI2BB2X1M U145 (.Y(n220), 
	.B1(n8), 
	.B0(FE_OFN5_n25), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][5] ));
   OAI2BB2X1M U146 (.Y(n222), 
	.B1(n9), 
	.B0(FE_OFN5_n25), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][5] ));
   OAI2BB2X1M U147 (.Y(n224), 
	.B1(n10), 
	.B0(FE_OFN5_n25), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][5] ));
   OAI2BB2X1M U148 (.Y(n226), 
	.B1(n11), 
	.B0(FE_OFN5_n25), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][5] ));
   OAI2BB2X1M U149 (.Y(n253), 
	.B1(n8), 
	.B0(FE_OFN6_n26), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][6] ));
   OAI2BB2X1M U150 (.Y(n255), 
	.B1(n9), 
	.B0(FE_OFN6_n26), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][6] ));
   OAI2BB2X1M U151 (.Y(n257), 
	.B1(n10), 
	.B0(FE_OFN6_n26), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][6] ));
   OAI2BB2X1M U152 (.Y(n259), 
	.B1(n11), 
	.B0(FE_OFN6_n26), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][6] ));
   OAI2BB2X1M U153 (.Y(n286), 
	.B1(n8), 
	.B0(FE_OFN7_n27), 
	.A1N(n8), 
	.A0N(\FIFO_MEM[4][7] ));
   OAI2BB2X1M U154 (.Y(n288), 
	.B1(n9), 
	.B0(FE_OFN7_n27), 
	.A1N(n9), 
	.A0N(\FIFO_MEM[5][7] ));
   OAI2BB2X1M U155 (.Y(n290), 
	.B1(n10), 
	.B0(FE_OFN7_n27), 
	.A1N(n10), 
	.A0N(\FIFO_MEM[6][7] ));
   OAI2BB2X1M U156 (.Y(n292), 
	.B1(n11), 
	.B0(FE_OFN7_n27), 
	.A1N(n11), 
	.A0N(\FIFO_MEM[7][7] ));
   OAI2BB2X1M U157 (.Y(n63), 
	.B1(n12), 
	.B0(FE_OFN0_n3), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][0] ));
   OAI2BB2X1M U158 (.Y(n71), 
	.B1(n16), 
	.B0(FE_OFN0_n3), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][0] ));
   OAI2BB2X1M U159 (.Y(n96), 
	.B1(n12), 
	.B0(FE_OFN1_n21), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][1] ));
   OAI2BB2X1M U160 (.Y(n104), 
	.B1(n16), 
	.B0(FE_OFN1_n21), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][1] ));
   OAI2BB2X1M U161 (.Y(n129), 
	.B1(n12), 
	.B0(FE_OFN2_n22), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][2] ));
   OAI2BB2X1M U162 (.Y(n137), 
	.B1(n16), 
	.B0(FE_OFN2_n22), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][2] ));
   OAI2BB2X1M U163 (.Y(n162), 
	.B1(n12), 
	.B0(FE_OFN3_n23), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][3] ));
   OAI2BB2X1M U164 (.Y(n170), 
	.B1(n16), 
	.B0(FE_OFN3_n23), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][3] ));
   OAI2BB2X1M U165 (.Y(n195), 
	.B1(n12), 
	.B0(FE_OFN4_n24), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][4] ));
   OAI2BB2X1M U166 (.Y(n203), 
	.B1(n16), 
	.B0(FE_OFN4_n24), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][4] ));
   OAI2BB2X1M U167 (.Y(n228), 
	.B1(n12), 
	.B0(FE_OFN5_n25), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][5] ));
   OAI2BB2X1M U168 (.Y(n236), 
	.B1(n16), 
	.B0(FE_OFN5_n25), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][5] ));
   OAI2BB2X1M U169 (.Y(n261), 
	.B1(n12), 
	.B0(FE_OFN6_n26), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][6] ));
   OAI2BB2X1M U170 (.Y(n269), 
	.B1(n16), 
	.B0(FE_OFN6_n26), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][6] ));
   OAI2BB2X1M U171 (.Y(n294), 
	.B1(n12), 
	.B0(FE_OFN7_n27), 
	.A1N(n12), 
	.A0N(\FIFO_MEM[8][7] ));
   OAI2BB2X1M U172 (.Y(n302), 
	.B1(n16), 
	.B0(FE_OFN7_n27), 
	.A1N(n16), 
	.A0N(\FIFO_MEM[12][7] ));
   OAI2BB2X1M U173 (.Y(n51), 
	.B1(n6), 
	.B0(FE_OFN0_n3), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][0] ));
   OAI2BB2X1M U174 (.Y(n53), 
	.B1(n7), 
	.B0(FE_OFN0_n3), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][0] ));
   OAI2BB2X1M U175 (.Y(n65), 
	.B1(n13), 
	.B0(FE_OFN0_n3), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][0] ));
   OAI2BB2X1M U320 (.Y(n73), 
	.B1(n17), 
	.B0(FE_OFN0_n3), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][0] ));
   OAI2BB2X1M U321 (.Y(n84), 
	.B1(n6), 
	.B0(FE_OFN1_n21), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][1] ));
   OAI2BB2X1M U322 (.Y(n86), 
	.B1(n7), 
	.B0(FE_OFN1_n21), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][1] ));
   OAI2BB2X1M U323 (.Y(n98), 
	.B1(n13), 
	.B0(FE_OFN1_n21), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][1] ));
   OAI2BB2X1M U324 (.Y(n106), 
	.B1(n17), 
	.B0(FE_OFN1_n21), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][1] ));
   OAI2BB2X1M U325 (.Y(n117), 
	.B1(n6), 
	.B0(FE_OFN2_n22), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][2] ));
   OAI2BB2X1M U326 (.Y(n119), 
	.B1(n7), 
	.B0(FE_OFN2_n22), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][2] ));
   OAI2BB2X1M U327 (.Y(n131), 
	.B1(n13), 
	.B0(FE_OFN2_n22), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][2] ));
   OAI2BB2X1M U328 (.Y(n139), 
	.B1(n17), 
	.B0(FE_OFN2_n22), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][2] ));
   OAI2BB2X1M U329 (.Y(n150), 
	.B1(n6), 
	.B0(FE_OFN3_n23), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][3] ));
   OAI2BB2X1M U330 (.Y(n152), 
	.B1(n7), 
	.B0(FE_OFN3_n23), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][3] ));
   OAI2BB2X1M U331 (.Y(n164), 
	.B1(n13), 
	.B0(FE_OFN3_n23), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][3] ));
   OAI2BB2X1M U332 (.Y(n172), 
	.B1(n17), 
	.B0(FE_OFN3_n23), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][3] ));
   OAI2BB2X1M U333 (.Y(n183), 
	.B1(n6), 
	.B0(FE_OFN4_n24), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][4] ));
   OAI2BB2X1M U334 (.Y(n185), 
	.B1(n7), 
	.B0(FE_OFN4_n24), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][4] ));
   OAI2BB2X1M U335 (.Y(n197), 
	.B1(n13), 
	.B0(FE_OFN4_n24), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][4] ));
   OAI2BB2X1M U336 (.Y(n205), 
	.B1(n17), 
	.B0(FE_OFN4_n24), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][4] ));
   OAI2BB2X1M U337 (.Y(n216), 
	.B1(n6), 
	.B0(FE_OFN5_n25), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][5] ));
   OAI2BB2X1M U338 (.Y(n218), 
	.B1(n7), 
	.B0(FE_OFN5_n25), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][5] ));
   OAI2BB2X1M U339 (.Y(n230), 
	.B1(n13), 
	.B0(FE_OFN5_n25), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][5] ));
   OAI2BB2X1M U340 (.Y(n238), 
	.B1(n17), 
	.B0(FE_OFN5_n25), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][5] ));
   OAI2BB2X1M U341 (.Y(n249), 
	.B1(n6), 
	.B0(FE_OFN6_n26), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][6] ));
   OAI2BB2X1M U342 (.Y(n251), 
	.B1(n7), 
	.B0(FE_OFN6_n26), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][6] ));
   OAI2BB2X1M U343 (.Y(n263), 
	.B1(n13), 
	.B0(FE_OFN6_n26), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][6] ));
   OAI2BB2X1M U344 (.Y(n271), 
	.B1(n17), 
	.B0(FE_OFN6_n26), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][6] ));
   OAI2BB2X1M U345 (.Y(n282), 
	.B1(n6), 
	.B0(FE_OFN7_n27), 
	.A1N(n6), 
	.A0N(\FIFO_MEM[2][7] ));
   OAI2BB2X1M U346 (.Y(n284), 
	.B1(n7), 
	.B0(FE_OFN7_n27), 
	.A1N(n7), 
	.A0N(\FIFO_MEM[3][7] ));
   OAI2BB2X1M U347 (.Y(n296), 
	.B1(n13), 
	.B0(FE_OFN7_n27), 
	.A1N(n13), 
	.A0N(\FIFO_MEM[9][7] ));
   OAI2BB2X1M U348 (.Y(n304), 
	.B1(n17), 
	.B0(FE_OFN7_n27), 
	.A1N(n17), 
	.A0N(\FIFO_MEM[13][7] ));
   OAI2BB2X1M U349 (.Y(n67), 
	.B1(n14), 
	.B0(FE_OFN0_n3), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][0] ));
   OAI2BB2X1M U350 (.Y(n69), 
	.B1(n15), 
	.B0(FE_OFN0_n3), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][0] ));
   OAI2BB2X1M U351 (.Y(n75), 
	.B1(n18), 
	.B0(FE_OFN0_n3), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][0] ));
   OAI2BB2X1M U352 (.Y(n77), 
	.B1(n19), 
	.B0(FE_OFN0_n3), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][0] ));
   OAI2BB2X1M U353 (.Y(n100), 
	.B1(n14), 
	.B0(FE_OFN1_n21), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][1] ));
   OAI2BB2X1M U354 (.Y(n102), 
	.B1(n15), 
	.B0(FE_OFN1_n21), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][1] ));
   OAI2BB2X1M U355 (.Y(n108), 
	.B1(n18), 
	.B0(FE_OFN1_n21), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][1] ));
   OAI2BB2X1M U356 (.Y(n110), 
	.B1(n19), 
	.B0(FE_OFN1_n21), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][1] ));
   OAI2BB2X1M U357 (.Y(n133), 
	.B1(n14), 
	.B0(FE_OFN2_n22), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][2] ));
   OAI2BB2X1M U358 (.Y(n135), 
	.B1(n15), 
	.B0(FE_OFN2_n22), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][2] ));
   OAI2BB2X1M U359 (.Y(n141), 
	.B1(n18), 
	.B0(FE_OFN2_n22), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][2] ));
   OAI2BB2X1M U360 (.Y(n143), 
	.B1(n19), 
	.B0(FE_OFN2_n22), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][2] ));
   OAI2BB2X1M U361 (.Y(n166), 
	.B1(n14), 
	.B0(FE_OFN3_n23), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][3] ));
   OAI2BB2X1M U362 (.Y(n168), 
	.B1(n15), 
	.B0(FE_OFN3_n23), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][3] ));
   OAI2BB2X1M U363 (.Y(n174), 
	.B1(n18), 
	.B0(FE_OFN3_n23), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][3] ));
   OAI2BB2X1M U364 (.Y(n176), 
	.B1(n19), 
	.B0(FE_OFN3_n23), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][3] ));
   OAI2BB2X1M U365 (.Y(n199), 
	.B1(n14), 
	.B0(FE_OFN4_n24), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][4] ));
   OAI2BB2X1M U366 (.Y(n201), 
	.B1(n15), 
	.B0(FE_OFN4_n24), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][4] ));
   OAI2BB2X1M U367 (.Y(n207), 
	.B1(n18), 
	.B0(FE_OFN4_n24), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][4] ));
   OAI2BB2X1M U368 (.Y(n209), 
	.B1(n19), 
	.B0(FE_OFN4_n24), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][4] ));
   OAI2BB2X1M U369 (.Y(n232), 
	.B1(n14), 
	.B0(FE_OFN5_n25), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][5] ));
   OAI2BB2X1M U370 (.Y(n234), 
	.B1(n15), 
	.B0(FE_OFN5_n25), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][5] ));
   OAI2BB2X1M U371 (.Y(n240), 
	.B1(n18), 
	.B0(FE_OFN5_n25), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][5] ));
   OAI2BB2X1M U372 (.Y(n242), 
	.B1(n19), 
	.B0(FE_OFN5_n25), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][5] ));
   OAI2BB2X1M U373 (.Y(n265), 
	.B1(n14), 
	.B0(FE_OFN6_n26), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][6] ));
   OAI2BB2X1M U374 (.Y(n267), 
	.B1(n15), 
	.B0(FE_OFN6_n26), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][6] ));
   OAI2BB2X1M U375 (.Y(n273), 
	.B1(n18), 
	.B0(FE_OFN6_n26), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][6] ));
   OAI2BB2X1M U376 (.Y(n275), 
	.B1(n19), 
	.B0(FE_OFN6_n26), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][6] ));
   OAI2BB2X1M U377 (.Y(n298), 
	.B1(n14), 
	.B0(FE_OFN7_n27), 
	.A1N(n14), 
	.A0N(\FIFO_MEM[10][7] ));
   OAI2BB2X1M U378 (.Y(n300), 
	.B1(n15), 
	.B0(FE_OFN7_n27), 
	.A1N(n15), 
	.A0N(\FIFO_MEM[11][7] ));
   OAI2BB2X1M U379 (.Y(n306), 
	.B1(n18), 
	.B0(FE_OFN7_n27), 
	.A1N(n18), 
	.A0N(\FIFO_MEM[14][7] ));
   OAI2BB2X1M U380 (.Y(n308), 
	.B1(n19), 
	.B0(FE_OFN7_n27), 
	.A1N(n19), 
	.A0N(\FIFO_MEM[15][7] ));
   MX4X1M U381 (.Y(n323), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[3][1] ), 
	.C(\FIFO_MEM[2][1] ), 
	.B(\FIFO_MEM[1][1] ), 
	.A(\FIFO_MEM[0][1] ));
   MX4X1M U382 (.Y(n318), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[7][0] ), 
	.C(\FIFO_MEM[6][0] ), 
	.B(\FIFO_MEM[5][0] ), 
	.A(\FIFO_MEM[4][0] ));
   MX4X1M U383 (.Y(n322), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[7][1] ), 
	.C(\FIFO_MEM[6][1] ), 
	.B(\FIFO_MEM[5][1] ), 
	.A(\FIFO_MEM[4][1] ));
   MX4X1M U384 (.Y(n326), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[7][2] ), 
	.C(\FIFO_MEM[6][2] ), 
	.B(\FIFO_MEM[5][2] ), 
	.A(\FIFO_MEM[4][2] ));
   MX4X1M U385 (.Y(n330), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[7][3] ), 
	.C(\FIFO_MEM[6][3] ), 
	.B(\FIFO_MEM[5][3] ), 
	.A(\FIFO_MEM[4][3] ));
   MX4X1M U386 (.Y(n334), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[7][4] ), 
	.C(\FIFO_MEM[6][4] ), 
	.B(\FIFO_MEM[5][4] ), 
	.A(\FIFO_MEM[4][4] ));
   MX4X1M U387 (.Y(n338), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[7][5] ), 
	.C(\FIFO_MEM[6][5] ), 
	.B(\FIFO_MEM[5][5] ), 
	.A(\FIFO_MEM[4][5] ));
   MX4X1M U388 (.Y(n342), 
	.S1(N12), 
	.S0(N11), 
	.D(\FIFO_MEM[7][6] ), 
	.C(\FIFO_MEM[6][6] ), 
	.B(\FIFO_MEM[5][6] ), 
	.A(\FIFO_MEM[4][6] ));
   MX4X1M U389 (.Y(n346), 
	.S1(N12), 
	.S0(n397), 
	.D(\FIFO_MEM[7][7] ), 
	.C(\FIFO_MEM[6][7] ), 
	.B(\FIFO_MEM[5][7] ), 
	.A(\FIFO_MEM[4][7] ));
   MX4X1M U390 (.Y(n360), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[7][1] ), 
	.C(\FIFO_MEM[6][1] ), 
	.B(\FIFO_MEM[5][1] ), 
	.A(\FIFO_MEM[4][1] ));
   MX4X1M U391 (.Y(n34), 
	.S1(n350), 
	.S0(N11), 
	.D(\FIFO_MEM[15][0] ), 
	.C(\FIFO_MEM[14][0] ), 
	.B(\FIFO_MEM[13][0] ), 
	.A(\FIFO_MEM[12][0] ));
   MX4X1M U392 (.Y(n354), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[15][0] ), 
	.C(\FIFO_MEM[14][0] ), 
	.B(\FIFO_MEM[13][0] ), 
	.A(\FIFO_MEM[12][0] ));
   MX4X1M U393 (.Y(n324), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[15][2] ), 
	.C(\FIFO_MEM[14][2] ), 
	.B(\FIFO_MEM[13][2] ), 
	.A(\FIFO_MEM[12][2] ));
   MX4X1M U394 (.Y(n328), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[15][3] ), 
	.C(\FIFO_MEM[14][3] ), 
	.B(\FIFO_MEM[13][3] ), 
	.A(\FIFO_MEM[12][3] ));
   MX4X1M U395 (.Y(n332), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[15][4] ), 
	.C(\FIFO_MEM[14][4] ), 
	.B(\FIFO_MEM[13][4] ), 
	.A(\FIFO_MEM[12][4] ));
   MX4X1M U396 (.Y(n336), 
	.S1(N12), 
	.S0(N11), 
	.D(\FIFO_MEM[15][5] ), 
	.C(\FIFO_MEM[14][5] ), 
	.B(\FIFO_MEM[13][5] ), 
	.A(\FIFO_MEM[12][5] ));
   MX4X1M U397 (.Y(n340), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[15][6] ), 
	.C(\FIFO_MEM[14][6] ), 
	.B(\FIFO_MEM[13][6] ), 
	.A(\FIFO_MEM[12][6] ));
   MX4X1M U398 (.Y(n344), 
	.S1(n350), 
	.S0(n397), 
	.D(\FIFO_MEM[15][7] ), 
	.C(\FIFO_MEM[14][7] ), 
	.B(\FIFO_MEM[13][7] ), 
	.A(\FIFO_MEM[12][7] ));
   MX4X1M U399 (.Y(n362), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[15][2] ), 
	.C(\FIFO_MEM[14][2] ), 
	.B(\FIFO_MEM[13][2] ), 
	.A(\FIFO_MEM[12][2] ));
   MX4X1M U400 (.Y(n366), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[15][3] ), 
	.C(\FIFO_MEM[14][3] ), 
	.B(\FIFO_MEM[13][3] ), 
	.A(\FIFO_MEM[12][3] ));
   MX4X1M U401 (.Y(n370), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[15][4] ), 
	.C(\FIFO_MEM[14][4] ), 
	.B(\FIFO_MEM[13][4] ), 
	.A(\FIFO_MEM[12][4] ));
   MX4X1M U402 (.Y(n374), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[15][5] ), 
	.C(\FIFO_MEM[14][5] ), 
	.B(\FIFO_MEM[13][5] ), 
	.A(\FIFO_MEM[12][5] ));
   MX4X1M U403 (.Y(n378), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[15][6] ), 
	.C(\FIFO_MEM[14][6] ), 
	.B(\FIFO_MEM[13][6] ), 
	.A(\FIFO_MEM[12][6] ));
   MX4X1M U404 (.Y(n382), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[15][7] ), 
	.C(\FIFO_MEM[14][7] ), 
	.B(\FIFO_MEM[13][7] ), 
	.A(\FIFO_MEM[12][7] ));
   MX4X1M U405 (.Y(N64), 
	.S1(N17), 
	.S0(N18), 
	.D(n354), 
	.C(n356), 
	.B(n355), 
	.A(n357));
   MX4X1M U406 (.Y(n357), 
	.S1(N16), 
	.S0(N15), 
	.D(\FIFO_MEM[3][0] ), 
	.C(\FIFO_MEM[2][0] ), 
	.B(\FIFO_MEM[1][0] ), 
	.A(\FIFO_MEM[0][0] ));
   MX4X1M U407 (.Y(n355), 
	.S1(N16), 
	.S0(N15), 
	.D(\FIFO_MEM[11][0] ), 
	.C(\FIFO_MEM[10][0] ), 
	.B(\FIFO_MEM[9][0] ), 
	.A(\FIFO_MEM[8][0] ));
   MX4X1M U408 (.Y(n356), 
	.S1(N16), 
	.S0(N15), 
	.D(\FIFO_MEM[7][0] ), 
	.C(\FIFO_MEM[6][0] ), 
	.B(\FIFO_MEM[5][0] ), 
	.A(\FIFO_MEM[4][0] ));
   MX4X1M U409 (.Y(N63), 
	.S1(N17), 
	.S0(N18), 
	.D(n358), 
	.C(n360), 
	.B(n359), 
	.A(n361));
   MX4X1M U410 (.Y(n359), 
	.S1(N16), 
	.S0(N15), 
	.D(\FIFO_MEM[11][1] ), 
	.C(\FIFO_MEM[10][1] ), 
	.B(\FIFO_MEM[9][1] ), 
	.A(\FIFO_MEM[8][1] ));
   MX4X1M U411 (.Y(n358), 
	.S1(n399), 
	.S0(n387), 
	.D(\FIFO_MEM[15][1] ), 
	.C(\FIFO_MEM[14][1] ), 
	.B(\FIFO_MEM[13][1] ), 
	.A(\FIFO_MEM[12][1] ));
   MX4X1M U412 (.Y(n361), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[3][1] ), 
	.C(\FIFO_MEM[2][1] ), 
	.B(\FIFO_MEM[1][1] ), 
	.A(\FIFO_MEM[0][1] ));
   MX4X1M U413 (.Y(N62), 
	.S1(N17), 
	.S0(N18), 
	.D(n362), 
	.C(n364), 
	.B(n363), 
	.A(n365));
   MX4X1M U414 (.Y(n365), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[3][2] ), 
	.C(\FIFO_MEM[2][2] ), 
	.B(\FIFO_MEM[1][2] ), 
	.A(\FIFO_MEM[0][2] ));
   MX4X1M U415 (.Y(n363), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[11][2] ), 
	.C(\FIFO_MEM[10][2] ), 
	.B(\FIFO_MEM[9][2] ), 
	.A(\FIFO_MEM[8][2] ));
   MX4X1M U416 (.Y(n364), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[7][2] ), 
	.C(\FIFO_MEM[6][2] ), 
	.B(\FIFO_MEM[5][2] ), 
	.A(\FIFO_MEM[4][2] ));
   MX4X1M U417 (.Y(N61), 
	.S1(N17), 
	.S0(N18), 
	.D(n366), 
	.C(n368), 
	.B(n367), 
	.A(n369));
   MX4X1M U418 (.Y(n369), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[3][3] ), 
	.C(\FIFO_MEM[2][3] ), 
	.B(\FIFO_MEM[1][3] ), 
	.A(\FIFO_MEM[0][3] ));
   MX4X1M U419 (.Y(n367), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[11][3] ), 
	.C(\FIFO_MEM[10][3] ), 
	.B(\FIFO_MEM[9][3] ), 
	.A(\FIFO_MEM[8][3] ));
   MX4X1M U420 (.Y(n368), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[7][3] ), 
	.C(\FIFO_MEM[6][3] ), 
	.B(\FIFO_MEM[5][3] ), 
	.A(\FIFO_MEM[4][3] ));
   MX4X1M U421 (.Y(N60), 
	.S1(N17), 
	.S0(N18), 
	.D(n370), 
	.C(n372), 
	.B(n371), 
	.A(n373));
   MX4X1M U422 (.Y(n373), 
	.S1(N16), 
	.S0(n388), 
	.D(\FIFO_MEM[3][4] ), 
	.C(\FIFO_MEM[2][4] ), 
	.B(\FIFO_MEM[1][4] ), 
	.A(\FIFO_MEM[0][4] ));
   MX4X1M U423 (.Y(n371), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[11][4] ), 
	.C(\FIFO_MEM[10][4] ), 
	.B(\FIFO_MEM[9][4] ), 
	.A(\FIFO_MEM[8][4] ));
   MX4X1M U424 (.Y(n372), 
	.S1(N16), 
	.S0(n387), 
	.D(\FIFO_MEM[7][4] ), 
	.C(\FIFO_MEM[6][4] ), 
	.B(\FIFO_MEM[5][4] ), 
	.A(\FIFO_MEM[4][4] ));
   MX4X1M U425 (.Y(N59), 
	.S1(N17), 
	.S0(N18), 
	.D(n374), 
	.C(n376), 
	.B(n375), 
	.A(n377));
   MX4X1M U426 (.Y(n377), 
	.S1(N16), 
	.S0(n388), 
	.D(\FIFO_MEM[3][5] ), 
	.C(\FIFO_MEM[2][5] ), 
	.B(\FIFO_MEM[1][5] ), 
	.A(\FIFO_MEM[0][5] ));
   MX4X1M U427 (.Y(n375), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[11][5] ), 
	.C(\FIFO_MEM[10][5] ), 
	.B(\FIFO_MEM[9][5] ), 
	.A(\FIFO_MEM[8][5] ));
   MX4X1M U428 (.Y(n376), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[7][5] ), 
	.C(\FIFO_MEM[6][5] ), 
	.B(\FIFO_MEM[5][5] ), 
	.A(\FIFO_MEM[4][5] ));
   MX4X1M U429 (.Y(N58), 
	.S1(N17), 
	.S0(N18), 
	.D(n378), 
	.C(n380), 
	.B(n379), 
	.A(n381));
   MX4X1M U430 (.Y(n381), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[3][6] ), 
	.C(\FIFO_MEM[2][6] ), 
	.B(\FIFO_MEM[1][6] ), 
	.A(\FIFO_MEM[0][6] ));
   MX4X1M U431 (.Y(n379), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[11][6] ), 
	.C(\FIFO_MEM[10][6] ), 
	.B(\FIFO_MEM[9][6] ), 
	.A(\FIFO_MEM[8][6] ));
   MX4X1M U432 (.Y(n380), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[7][6] ), 
	.C(\FIFO_MEM[6][6] ), 
	.B(\FIFO_MEM[5][6] ), 
	.A(\FIFO_MEM[4][6] ));
   MX4X1M U433 (.Y(N57), 
	.S1(N17), 
	.S0(N18), 
	.D(n382), 
	.C(n384), 
	.B(n383), 
	.A(n385));
   MX4X1M U434 (.Y(n385), 
	.S1(N16), 
	.S0(n388), 
	.D(\FIFO_MEM[3][7] ), 
	.C(\FIFO_MEM[2][7] ), 
	.B(\FIFO_MEM[1][7] ), 
	.A(\FIFO_MEM[0][7] ));
   MX4X1M U435 (.Y(n383), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[11][7] ), 
	.C(\FIFO_MEM[10][7] ), 
	.B(\FIFO_MEM[9][7] ), 
	.A(\FIFO_MEM[8][7] ));
   MX4X1M U436 (.Y(n384), 
	.S1(n399), 
	.S0(n388), 
	.D(\FIFO_MEM[7][7] ), 
	.C(\FIFO_MEM[6][7] ), 
	.B(\FIFO_MEM[5][7] ), 
	.A(\FIFO_MEM[4][7] ));
   INVX2M U437 (.Y(n399), 
	.A(n400));
   INVX2M U438 (.Y(n400), 
	.A(N16));
endmodule

module ASYNC_FIFO_test_1 (
	W_CLK, 
	W_RST, 
	W_INC, 
	R_CLK, 
	R_RST, 
	R_INC, 
	WR_DATA, 
	FULL, 
	EMPTY, 
	RD_DATA, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so3, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN10_RST_D1_M, 
	FE_OFN11_RST_D1_M, 
	FE_OFN12_RST_D1_M, 
	FE_OFN17_SE, 
	FE_OFN18_SE, 
	FE_OFN21_SE, 
	FE_OFN24_SE, 
	REF_CLK_M__L5_N2, 
	REF_CLK_M__L5_N3, 
	REF_CLK_M__L5_N4, 
	REF_CLK_M__L5_N7);
   input W_CLK;
   input W_RST;
   input W_INC;
   input R_CLK;
   input R_RST;
   input R_INC;
   input [7:0] WR_DATA;
   output FULL;
   output EMPTY;
   output [7:0] RD_DATA;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so3;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN10_RST_D1_M;
   input FE_OFN11_RST_D1_M;
   input FE_OFN12_RST_D1_M;
   input FE_OFN17_SE;
   input FE_OFN18_SE;
   input FE_OFN21_SE;
   input FE_OFN24_SE;
   input REF_CLK_M__L5_N2;
   input REF_CLK_M__L5_N3;
   input REF_CLK_M__L5_N4;
   input REF_CLK_M__L5_N7;

   // Internal wires
   wire wclk_en;
   wire rclk_en;
   wire n1;
   wire n2;
   wire n7;
   wire n8;
   wire n11;
   wire n12;
   wire [4:0] Wptr;
   wire [4:0] Wptr_sync;
   wire [4:0] Rptr;
   wire [4:0] Rptr_sync;
   wire [3:0] Waddr;
   wire [3:0] raddr;
   wire SYNOPSYS_UNCONNECTED__0;
   wire SYNOPSYS_UNCONNECTED__1;

   AND3X2M U2 (.Y(wclk_en), 
	.C(FE_OFN12_RST_D1_M), 
	.B(W_INC), 
	.A(n7));
   INVX2M U3 (.Y(n7), 
	.A(FULL));
   BUFX2M U4 (.Y(n1), 
	.A(Waddr[0]));
   AND3X2M U9 (.Y(rclk_en), 
	.C(R_RST), 
	.B(R_INC), 
	.A(n8));
   INVXLM U10 (.Y(n8), 
	.A(EMPTY));
   BUFX4M U11 (.Y(n2), 
	.A(Waddr[1]));
   Bit_Sync_00000002_00000005_test_1 sync_w2r (.RST_n(R_RST), 
	.CLK(R_CLK), 
	.ASYNC({ 1'b0,
		Wptr[3],
		Wptr[2],
		Wptr[1],
		Wptr[0] }), 
	.SYNC({ Wptr_sync[4],
		Wptr_sync[3],
		Wptr_sync[2],
		Wptr_sync[1],
		Wptr_sync[0] }), 
	.test_si2(test_si3), 
	.test_si1(n11), 
	.test_so2(test_so3), 
	.test_so1(test_so2), 
	.test_se(FE_OFN17_SE), 
	.FE_OFN18_SE(FE_OFN18_SE));
   Bit_Sync_00000002_00000005_test_0 sync_r2w (.RST_n(FE_OFN10_RST_D1_M), 
	.CLK(W_CLK), 
	.ASYNC({ 1'b0,
		Rptr[3],
		Rptr[2],
		Rptr[1],
		Rptr[0] }), 
	.SYNC({ Rptr_sync[4],
		Rptr_sync[3],
		Rptr_sync[2],
		Rptr_sync[1],
		Rptr_sync[0] }), 
	.test_si(Wptr[3]), 
	.test_so(n11), 
	.test_se(test_se), 
	.FE_OFN17_SE(FE_OFN17_SE), 
	.FE_OFN18_SE(FE_OFN18_SE));
   fifo_wrptr_full_00000008_00000010_test_1 fifo_wrptr_full_dut (.W_CLK(W_CLK), 
	.W_RST(FE_OFN10_RST_D1_M), 
	.W_INC(W_INC), 
	.gray_Rptr({ Rptr_sync[4],
		Rptr_sync[3],
		Rptr_sync[2],
		Rptr_sync[1],
		Rptr_sync[0] }), 
	.WFULL(FULL), 
	.Waddr({ Waddr[3],
		Waddr[2],
		Waddr[1],
		Waddr[0] }), 
	.gray_Wptr({ SYNOPSYS_UNCONNECTED__0,
		Wptr[3],
		Wptr[2],
		Wptr[1],
		Wptr[0] }), 
	.test_si(Rptr[3]), 
	.test_se(test_se), 
	.FE_OFN11_RST_D1_M(FE_OFN11_RST_D1_M), 
	.FE_OFN12_RST_D1_M(FE_OFN12_RST_D1_M), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.FE_OFN21_SE(FE_OFN21_SE), 
	.REF_CLK_M__L5_N2(REF_CLK_M__L5_N2));
   fifo_rdptr_empty_00000008_00000010_test_1 fifo_rdptr_empty_dut (.R_CLK(R_CLK), 
	.R_RST(R_RST), 
	.R_INC(R_INC), 
	.gray_Wptr({ Wptr_sync[4],
		Wptr_sync[3],
		Wptr_sync[2],
		Wptr_sync[1],
		Wptr_sync[0] }), 
	.REMPTY(EMPTY), 
	.Raddr({ raddr[3],
		raddr[2],
		raddr[1],
		raddr[0] }), 
	.gray_Rptr({ SYNOPSYS_UNCONNECTED__1,
		Rptr[3],
		Rptr[2],
		Rptr[1],
		Rptr[0] }), 
	.test_si(n12), 
	.test_se(FE_OFN17_SE), 
	.FE_OFN18_SE(FE_OFN18_SE), 
	.FE_OFN24_SE(FE_OFN24_SE));
   FIFO_MEMORY_00000008_00000010_test_1 FIFO_MEMORY_dut (.WCLK(W_CLK), 
	.WRST(W_RST), 
	.R_CLK(R_CLK), 
	.R_RST(R_RST), 
	.wdata({ WR_DATA[7],
		WR_DATA[6],
		WR_DATA[5],
		WR_DATA[4],
		WR_DATA[3],
		WR_DATA[2],
		WR_DATA[1],
		WR_DATA[0] }), 
	.wclk_en(wclk_en), 
	.rclk_en(rclk_en), 
	.waddr({ Waddr[3],
		Waddr[2],
		n2,
		n1 }), 
	.raddr({ raddr[3],
		raddr[2],
		raddr[1],
		raddr[0] }), 
	.rdata({ RD_DATA[7],
		RD_DATA[6],
		RD_DATA[5],
		RD_DATA[4],
		RD_DATA[3],
		RD_DATA[2],
		RD_DATA[1],
		RD_DATA[0] }), 
	.test_si2(test_si2), 
	.test_si1(test_si1), 
	.test_so2(n12), 
	.test_so1(test_so1), 
	.test_se(test_se), 
	.FE_OFN11_RST_D1_M(FE_OFN11_RST_D1_M), 
	.FE_OFN12_RST_D1_M(FE_OFN12_RST_D1_M), 
	.FE_OFN17_SE(FE_OFN17_SE), 
	.FE_OFN21_SE(FE_OFN21_SE), 
	.FE_OFN24_SE(FE_OFN24_SE), 
	.REF_CLK_M__L5_N2(REF_CLK_M__L5_N2), 
	.REF_CLK_M__L5_N3(REF_CLK_M__L5_N3), 
	.REF_CLK_M__L5_N4(REF_CLK_M__L5_N4), 
	.REF_CLK_M__L5_N7(REF_CLK_M__L5_N7));
endmodule

module PULSE_GENERATOR_test_1 (
	CLK, 
	RST_n, 
	in, 
	out, 
	test_si, 
	test_se);
   input CLK;
   input RST_n;
   input in;
   output out;
   input test_si;
   input test_se;

   // Internal wires
   wire Q_in;
   wire N1;

   SDFFRQX2M Q_in_reg (.SI(test_si), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(Q_in), 
	.D(in), 
	.CK(CLK));
   SDFFRQX2M out_reg (.SI(Q_in), 
	.SE(test_se), 
	.RN(RST_n), 
	.Q(out), 
	.D(N1), 
	.CK(CLK));
   NOR2BX2M U5 (.Y(N1), 
	.B(Q_in), 
	.AN(in));
endmodule

