`timescale 1ns / 1fs                     // 1ns -- 1000000 precision (6 numbers prescision)


module SYS_TOP_tb();


 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
 ///////////////////////////////////////////////////// PARAMETERS ///////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



 parameter REF_CLK_PERIOD  =  10           ;        //100MHZ
 parameter UART_CLK_PERIOD =  271.2673611  ;        // 3.6864 MHZ  , FOR PRESCALE = 1 -> 271.2673611 , PRESCALE = 2 -> 135.6336806
 parameter RX_CLK_PERIOD   =  135.6336806  ;        // 115.200 KHZ
 parameter TX_CLK_PERIOD   =  8680.555556  ;
 
 parameter PRESCALE = 'd16                 ;



 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
 ////////////////////////////////////////////// CONEECTIONS DECLARATION /////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

 reg REF_CLK     ;
 reg UART_CLK    ;
 reg RST         ;
 reg RX_IN       ;

 wire TX_OUT     ;

 wire RX_CLK     ;
 wire TX_CLK     ;

 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
 ////////////////////////////////////////////////// STIMULUS MEMORY /////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


reg Data_Seed_Write_RF_h           [32:0];
reg Data_Seed_Write_ALU_CMD_h      [43:0];
reg Data_Seed_Read_RF_h            [21:0];
reg Data_Seed_Write_ALU_No_CMD_h   [21:0];


 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
 ////////////////////////////////////////////// CONEECTIONS DECLARATION /////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


integer i ;
integer j ;
integer k ;
integer n ;
 

 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
 ////////////////////////////////////////////// TOP_MODULE INSTANTIATION ////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 //////////////////////////////////////////////////////////////////////////////////////////////////////////////////////// 



SYS_TOP SYS_TOP_dut
(
 .REF_CLK  (REF_CLK)     ,
 .UART_CLK (UART_CLK)    ,
 .RST      (RST)         ,
 .RX_IN    (RX_IN)       ,

 .TX_OUT   (TX_OUT)
);



 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
 ////////////////////////////////////////////// CLOCK DOMAINS GENERATION ////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 //////////////////////////////////////////////////////////////////////////////////////////////////////////////////////// 


  always begin
    #(REF_CLK_PERIOD / 2)   REF_CLK  = ~ REF_CLK   ;
  end



  always begin
    #(UART_CLK_PERIOD / 2)  UART_CLK = ~ UART_CLK  ;
  end


 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////	
 ////////////////////////////////////////////// CLOCK DOMAINS GENERATION ////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



ClkDiv__ CLK_DIV_RX_dut
(
.i_ref_clk   (UART_CLK),
.i_rst_n     (RST_D2),
.i_div_ratio (2),

.o_div_clk(RX_CLK)
);


ClkDiv__ CLK_DIV_TX_dut
(
.i_ref_clk   (UART_CLK),
.i_rst_n     (RST_D2),
.i_div_ratio (32),

.o_div_clk(TX_CLK)
);





Rst_Sync #(.NUM_STAGES(2) , .ACTIVE_TYP("LOW")) Rst_Sync_D1_dut (

.RST       (RST),
.CLK       (REF_CLK),
.SYNC_RST  (RST_D1)

);



Rst_Sync #(.NUM_STAGES(2) , .ACTIVE_TYP("LOW")) Rst_Sync_D2_dut (

.RST       (RST),
.CLK       (UART_CLK),
.SYNC_RST  (RST_D2)

);









///////////////////////////////////////////////////


 initial begin

     $readmemh ("Data_Seed_Write_RF_h.txt" , Data_Seed_Write_RF_h );
     $readmemh("Data_Seed_Write_ALU_CMD_h.txt",Data_Seed_Write_ALU_CMD_h);
     $readmemh("Data_Seed_Read_RF_h.txt", Data_Seed_Read_RF_h);
     $readmemh("Data_Seed_Write_ALU_No_CMD_h.txt",Data_Seed_Write_ALU_No_CMD_h);
   
    // Initialize inputs
    REF_CLK = 0;
    UART_CLK =0;
    RX_IN = 0;
    i = 0 ;
    j = 0;
    k = 0; 
    n =0 ;
    
    // R_INC = 0 ;
    // bus_enable = 0;
    // data_in_syn = 8'h00;
    //enable_pulse = 0;
    // FIFO_FULL = 0;
    // // Rd_DATA = 8'h00;
    // Rd_Valid = 0;
    // ALU_OUT = 16'h0000;
    // OUT_VALID = 0;
     
     RST = 0; 
    // Release reset
    #(REF_CLK_PERIOD) RST = 1; 
    #(2*REF_CLK_PERIOD);
    




//=============== WRITE IN RF =========================


      for(i = 0 ; i < 11 ; i = i + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_RF_h[i];
      repeat(PRESCALE) @(negedge RX_CLK);
      end


      #(RX_CLK_PERIOD) ;


      for(i = 11 ; i < 22 ; i = i + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_RF_h[i];
      repeat(PRESCALE) @(negedge RX_CLK);
      end

     #(RX_CLK_PERIOD) ;

    
      for(i = 22 ; i < 33 ; i = i + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_RF_h[i];
      repeat(PRESCALE) @(negedge RX_CLK);
      end
      
      
      #(RX_CLK_PERIOD) ;


       
  //=================================================



//=============== WRITE IN ALU WITH CMD ================


      for(j = 0 ; j < 11 ; j = j + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_ALU_CMD_h[j];
      repeat(PRESCALE) @(negedge RX_CLK);
      end


      #(RX_CLK_PERIOD) ;


      for(j = 11 ; j < 22 ; j = j + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_ALU_CMD_h[j];
      repeat(PRESCALE) @(negedge RX_CLK);
      end

     #(RX_CLK_PERIOD) ;

    
      for(j = 22 ; j < 33 ; j = j + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_ALU_CMD_h[j];
      repeat(PRESCALE) @(negedge RX_CLK);
      end
      
      
      #(RX_CLK_PERIOD) ;



      for(j = 33 ; j < 44 ; j = j + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_ALU_CMD_h[j];
      repeat(PRESCALE) @(negedge RX_CLK);
      end
      
      
      #(RX_CLK_PERIOD) ;


       
  //====================================================


  //=============== READ FROM RF ===============

   
      for(k = 0 ; k < 11 ; k = k + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Read_RF_h[k];
      repeat(PRESCALE) @(negedge RX_CLK);
      end
      
      
      #(RX_CLK_PERIOD) ;



      for(k = 11 ; k < 22 ; k = k + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Read_RF_h[k];
      repeat(PRESCALE) @(negedge RX_CLK);
      end
      
      
      #(RX_CLK_PERIOD) ;
   

  //============================================

  //=======  WRITE IN ALU WITH No OPERAND ======

   
      for(n = 0 ; n < 11 ; n = n + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_ALU_No_CMD_h[n];
      repeat(PRESCALE) @(negedge RX_CLK);
      end
      
      
      #(RX_CLK_PERIOD) ;


      for(n = 11 ; n < 22 ; n = n + 1)
      begin
      @(negedge RX_CLK);
      RX_IN = Data_Seed_Write_ALU_No_CMD_h[n];
      repeat(PRESCALE) @(negedge RX_CLK);
      end
      
      
      #(RX_CLK_PERIOD) ;

      
      // R_INC = 1'b1;

       #(20*TX_CLK_PERIOD);

      // R_INC = 0;

    //  RST = 0; 
    // // Release reset
    // //#(REF_CLK_PERIOD) RST = 1; 
    // #(2*REF_CLK_PERIOD);

  //============================================
      


    #50 $stop;
  end




////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////// CLOCK DOMAINS GENERATION ////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


task initialize();
 begin	

    REF_CLK  = 0 ;
    UART_CLK = 0 ;
    RX_IN    = 0 ;

 end	
endtask 



task RESET();
 begin
 	
    RST = 0 ;
    #(2*REF_CLK_PERIOD) ; 
    RST = 1 ; 
    #(2*REF_CLK_PERIOD) ;

 end
endtask 



task transmit(input Data_in);
 begin
 	
 	RX_IN = Data_in ;
 	// repeat(PRESCALE) @(negedge rst_n);


 end
endtask




endmodule